magic
tech sky130A
magscale 1 2
timestamp 1746986264
<< obsli1 >>
rect -1580 7722 1730 7804
rect -1580 -1722 -1498 7722
rect -798 6757 948 7022
rect -798 -757 -716 6757
rect -659 -164 -457 6165
rect -134 -164 284 6165
rect 607 -164 809 6165
rect -146 -657 290 -443
rect 866 -757 948 6757
rect -798 -1022 948 -757
rect 1648 -1722 1730 7722
rect -1580 -1804 1730 -1722
<< obsm1 >>
rect -1580 7722 1730 7804
rect -1580 -1722 -1498 7722
rect -798 6757 948 7022
rect -798 -757 -716 6757
rect -659 -164 -457 6165
rect -134 -164 284 6165
rect 607 -164 809 6165
rect -146 -657 290 -443
rect 866 -757 948 6757
rect -798 -1022 948 -757
rect 1648 -1722 1730 7722
rect -1580 -1804 1730 -1722
<< obsm2 >>
rect -659 -1122 -457 6165
rect -134 -164 284 7122
rect -146 -657 290 -443
rect 607 -1122 809 6165
<< obsm3 >>
rect -150 -657 290 -443
<< properties >>
string FIXED_BBOX 0 0 3310 9608
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10317996
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10046666
<< end >>
