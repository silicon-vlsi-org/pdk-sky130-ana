magic
tech sky130A
magscale 1 2
timestamp 1746986264
<< locali >>
rect 191 752 195 786
rect 229 752 267 786
rect 301 752 339 786
rect 373 752 411 786
rect 445 752 483 786
rect 517 752 555 786
rect 589 752 627 786
rect 661 752 665 786
rect 48 672 82 674
rect 48 600 82 638
rect 48 528 82 566
rect 48 456 82 494
rect 48 384 82 422
rect 48 312 82 350
rect 48 240 82 278
rect 48 168 82 206
rect 48 132 82 134
rect 774 672 808 674
rect 774 600 808 638
rect 774 528 808 566
rect 774 456 808 494
rect 774 384 808 422
rect 774 312 808 350
rect 774 240 808 278
rect 774 168 808 206
rect 774 132 808 134
rect 191 20 195 54
rect 229 20 267 54
rect 301 20 339 54
rect 373 20 411 54
rect 445 20 483 54
rect 517 20 555 54
rect 589 20 627 54
rect 661 20 665 54
<< viali >>
rect 195 752 229 786
rect 267 752 301 786
rect 339 752 373 786
rect 411 752 445 786
rect 483 752 517 786
rect 555 752 589 786
rect 627 752 661 786
rect 48 638 82 672
rect 48 566 82 600
rect 48 494 82 528
rect 48 422 82 456
rect 48 350 82 384
rect 48 278 82 312
rect 48 206 82 240
rect 48 134 82 168
rect 774 638 808 672
rect 774 566 808 600
rect 774 494 808 528
rect 774 422 808 456
rect 774 350 808 384
rect 774 278 808 312
rect 774 206 808 240
rect 774 134 808 168
rect 195 20 229 54
rect 267 20 301 54
rect 339 20 373 54
rect 411 20 445 54
rect 483 20 517 54
rect 555 20 589 54
rect 627 20 661 54
<< obsli1 >>
rect 159 98 193 708
rect 285 98 319 708
rect 411 98 445 708
rect 537 98 571 708
rect 663 98 697 708
<< metal1 >>
rect 183 786 673 806
rect 183 752 195 786
rect 229 752 267 786
rect 301 752 339 786
rect 373 752 411 786
rect 445 752 483 786
rect 517 752 555 786
rect 589 752 627 786
rect 661 752 673 786
rect 183 740 673 752
rect 36 672 94 684
rect 36 638 48 672
rect 82 638 94 672
rect 36 600 94 638
rect 36 566 48 600
rect 82 566 94 600
rect 36 528 94 566
rect 36 494 48 528
rect 82 494 94 528
rect 36 456 94 494
rect 36 422 48 456
rect 82 422 94 456
rect 36 384 94 422
rect 36 350 48 384
rect 82 350 94 384
rect 36 312 94 350
rect 36 278 48 312
rect 82 278 94 312
rect 36 240 94 278
rect 36 206 48 240
rect 82 206 94 240
rect 36 168 94 206
rect 36 134 48 168
rect 82 134 94 168
rect 36 122 94 134
rect 762 672 820 684
rect 762 638 774 672
rect 808 638 820 672
rect 762 600 820 638
rect 762 566 774 600
rect 808 566 820 600
rect 762 528 820 566
rect 762 494 774 528
rect 808 494 820 528
rect 762 456 820 494
rect 762 422 774 456
rect 808 422 820 456
rect 762 384 820 422
rect 762 350 774 384
rect 808 350 820 384
rect 762 312 820 350
rect 762 278 774 312
rect 808 278 820 312
rect 762 240 820 278
rect 762 206 774 240
rect 808 206 820 240
rect 762 168 820 206
rect 762 134 774 168
rect 808 134 820 168
rect 762 122 820 134
rect 183 54 673 66
rect 183 20 195 54
rect 229 20 267 54
rect 301 20 339 54
rect 373 20 411 54
rect 445 20 483 54
rect 517 20 555 54
rect 589 20 627 54
rect 661 20 673 54
rect 183 0 673 20
<< obsm1 >>
rect 150 122 202 684
rect 276 122 328 684
rect 402 122 454 684
rect 528 122 580 684
rect 654 122 706 684
<< metal2 >>
rect 10 428 846 684
rect 10 122 846 378
<< labels >>
rlabel viali s 774 638 808 672 6 BULK
port 1 nsew
rlabel viali s 774 566 808 600 6 BULK
port 1 nsew
rlabel viali s 774 494 808 528 6 BULK
port 1 nsew
rlabel viali s 774 422 808 456 6 BULK
port 1 nsew
rlabel viali s 774 350 808 384 6 BULK
port 1 nsew
rlabel viali s 774 278 808 312 6 BULK
port 1 nsew
rlabel viali s 774 206 808 240 6 BULK
port 1 nsew
rlabel viali s 774 134 808 168 6 BULK
port 1 nsew
rlabel viali s 48 638 82 672 6 BULK
port 1 nsew
rlabel viali s 48 566 82 600 6 BULK
port 1 nsew
rlabel viali s 48 494 82 528 6 BULK
port 1 nsew
rlabel viali s 48 422 82 456 6 BULK
port 1 nsew
rlabel viali s 48 350 82 384 6 BULK
port 1 nsew
rlabel viali s 48 278 82 312 6 BULK
port 1 nsew
rlabel viali s 48 206 82 240 6 BULK
port 1 nsew
rlabel viali s 48 134 82 168 6 BULK
port 1 nsew
rlabel locali s 774 132 808 674 6 BULK
port 1 nsew
rlabel locali s 48 132 82 674 6 BULK
port 1 nsew
rlabel metal1 s 762 122 820 684 6 BULK
port 1 nsew
rlabel metal1 s 36 122 94 684 6 BULK
port 1 nsew
rlabel metal2 s 10 428 846 684 6 DRAIN
port 2 nsew
rlabel viali s 627 752 661 786 6 GATE
port 3 nsew
rlabel viali s 627 20 661 54 6 GATE
port 3 nsew
rlabel viali s 555 752 589 786 6 GATE
port 3 nsew
rlabel viali s 555 20 589 54 6 GATE
port 3 nsew
rlabel viali s 483 752 517 786 6 GATE
port 3 nsew
rlabel viali s 483 20 517 54 6 GATE
port 3 nsew
rlabel viali s 411 752 445 786 6 GATE
port 3 nsew
rlabel viali s 411 20 445 54 6 GATE
port 3 nsew
rlabel viali s 339 752 373 786 6 GATE
port 3 nsew
rlabel viali s 339 20 373 54 6 GATE
port 3 nsew
rlabel viali s 267 752 301 786 6 GATE
port 3 nsew
rlabel viali s 267 20 301 54 6 GATE
port 3 nsew
rlabel viali s 195 752 229 786 6 GATE
port 3 nsew
rlabel viali s 195 20 229 54 6 GATE
port 3 nsew
rlabel locali s 191 752 665 786 6 GATE
port 3 nsew
rlabel locali s 191 20 665 54 6 GATE
port 3 nsew
rlabel metal1 s 183 740 673 806 6 GATE
port 3 nsew
rlabel metal1 s 183 0 673 66 6 GATE
port 3 nsew
rlabel metal2 s 10 122 846 378 6 SOURCE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 856 806
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9931810
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9916306
<< end >>
