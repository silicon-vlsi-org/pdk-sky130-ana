* SKY130 Spice File.
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__special_nfet_01v8__ff.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__special_nfet_01v8__mismatch.corner.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__special_pfet_01v8_hvt__ff.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__special_pfet_01v8_hvt__mismatch.corner.spice"
.include "all.spice"
.include "ff/legacy.spice"
.include "ff/nonfet.spice"
.include "ff/rf.spice"
