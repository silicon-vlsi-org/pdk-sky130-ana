magic
tech sky130A
magscale 1 2
timestamp 1746986264
<< obsm2 >>
rect -7432 31006 -987 33506
tri -987 31006 1513 33506 sw
tri -2023 28004 979 31006 ne
rect 979 30504 1513 31006
tri 1513 30504 2015 31006 sw
rect 979 28004 7787 30504
rect -7432 25002 -987 27502
tri -987 25002 1513 27502 sw
tri -2023 22000 979 25002 ne
rect 979 24500 1513 25002
tri 1513 24500 2015 25002 sw
rect 979 22000 7787 24500
rect 19408 -1250 37508 1250
tri -2023 -28004 979 -25002 se
rect 979 -27502 7675 -25002
rect 979 -28004 1513 -27502
tri 1513 -28004 2015 -27502 nw
rect -7544 -30504 -987 -28004
tri -987 -30504 1513 -28004 nw
tri -2023 -34008 979 -31006 se
rect 979 -33506 7675 -31006
rect 979 -34008 1513 -33506
tri 1513 -34008 2015 -33506 nw
rect -7544 -36508 -987 -34008
tri -987 -36508 1513 -34008 nw
<< obsm3 >>
tri -17624 34008 -15124 36508 se
rect -15124 34008 15124 36508
tri 15124 34008 17624 36508 sw
tri -20305 31327 -17624 34008 se
rect -17624 33506 -14590 34008
tri -14590 33506 -14088 34008 nw
tri 14088 33506 14590 34008 ne
rect 14590 33506 17624 34008
rect -17624 32804 -15292 33506
tri -15292 32804 -14590 33506 nw
tri -14583 32804 -13881 33506 se
rect -13881 33286 -2268 33506
tri -2268 33286 -2048 33506 sw
rect -13881 32804 -2048 33286
tri 285 32804 987 33506 se
rect 987 32804 13881 33506
tri 13881 32804 14583 33506 sw
tri 14590 32804 15292 33506 ne
rect 15292 32804 17624 33506
rect -17624 32095 -16001 32804
tri -16001 32095 -15292 32804 nw
tri -15292 32095 -14583 32804 se
rect -14583 32095 -2048 32804
rect -17624 31388 -16708 32095
tri -16708 31388 -16001 32095 nw
tri -15999 31388 -15292 32095 se
rect -15292 31388 -2048 32095
rect -17624 31327 -17417 31388
tri -23307 28325 -20305 31327 se
rect -20305 30679 -17417 31327
tri -17417 30679 -16708 31388 nw
tri -16708 30679 -15999 31388 se
rect -15999 31226 -2048 31388
rect -15999 31006 -2268 31226
tri -2268 31006 -2048 31226 nw
rect -15999 30679 -13534 31006
rect -20305 29970 -18126 30679
tri -18126 29970 -17417 30679 nw
tri -17417 29970 -16708 30679 se
rect -16708 30317 -13534 30679
tri -13534 30317 -12845 31006 nw
tri -2015 30504 285 32804 se
rect 285 32270 14583 32804
tri 14583 32270 15117 32804 sw
tri 15292 32270 15826 32804 ne
rect 15826 32270 17624 32804
rect 285 31561 15117 32270
tri 15117 31561 15826 32270 sw
tri 15826 31561 16535 32270 ne
rect 16535 31561 17624 32270
tri 17624 31561 20071 34008 sw
rect 285 31006 15826 31561
tri -12824 30317 -12637 30504 se
rect -12637 30317 285 30504
rect -16708 29970 -14162 30317
rect -20305 29268 -18828 29970
tri -18828 29268 -18126 29970 nw
tri -18119 29268 -17417 29970 se
rect -17417 29689 -14162 29970
tri -14162 29689 -13534 30317 nw
tri -13452 29689 -12824 30317 se
rect -12824 29689 285 30317
rect -17417 29268 -14776 29689
rect -20305 28559 -19537 29268
tri -19537 28559 -18828 29268 nw
tri -18828 28559 -18119 29268 se
rect -18119 29075 -14776 29268
tri -14776 29075 -14162 29689 nw
tri -14066 29075 -13452 29689 se
rect -13452 29268 285 29689
tri 285 29268 2023 31006 nw
tri 12845 30504 13347 31006 ne
rect 13347 30852 15826 31006
tri 15826 30852 16535 31561 sw
tri 16535 30852 17244 31561 ne
rect 17244 30852 20071 31561
rect 13347 30504 16535 30852
tri 2403 30284 2623 30504 se
rect 2623 30284 12637 30504
rect 2403 29970 12637 30284
tri 12637 29970 13171 30504 sw
tri 13347 29970 13881 30504 ne
rect 13881 30143 16535 30504
tri 16535 30143 17244 30852 sw
tri 17244 30143 17953 30852 ne
rect 17953 30143 20071 30852
rect 13881 29970 17244 30143
rect 2403 29268 13171 29970
tri 13171 29268 13873 29970 sw
tri 13881 29268 14583 29970 ne
rect 14583 29436 17244 29970
tri 17244 29436 17951 30143 sw
tri 17953 29436 18660 30143 ne
rect 18660 29436 20071 30143
rect 14583 29268 17951 29436
rect -13452 29075 -979 29268
rect -18119 28559 -15293 29075
rect -20305 28325 -20244 28559
tri -26309 25323 -23307 28325 se
rect -23307 27852 -20244 28325
tri -20244 27852 -19537 28559 nw
tri -19535 27852 -18828 28559 se
rect -18828 28558 -15293 28559
tri -15293 28558 -14776 29075 nw
tri -14583 28558 -14066 29075 se
rect -14066 28558 -979 29075
rect -18828 28025 -15826 28558
tri -15826 28025 -15293 28558 nw
tri -15116 28025 -14583 28558 se
rect -14583 28025 -979 28558
rect -18828 27852 -16173 28025
rect -23307 27143 -20953 27852
tri -20953 27143 -20244 27852 nw
tri -20244 27143 -19535 27852 se
rect -19535 27678 -16173 27852
tri -16173 27678 -15826 28025 nw
tri -15463 27678 -15116 28025 se
rect -15116 28004 -979 28025
tri -979 28004 285 29268 nw
rect 2403 28558 13873 29268
tri 13873 28558 14583 29268 sw
tri 14583 28558 15293 29268 ne
rect 15293 28734 17951 29268
tri 17951 28734 18653 29436 sw
tri 18660 28734 19362 29436 ne
rect 19362 28734 20071 29436
rect 15293 28558 18653 28734
rect 2403 28224 14583 28558
tri 2403 28004 2623 28224 ne
rect 2623 28025 14583 28224
tri 14583 28025 15116 28558 sw
tri 15293 28025 15826 28558 ne
rect 15826 28025 18653 28558
tri 18653 28025 19362 28734 sw
tri 19362 28025 20071 28734 ne
tri 20071 28025 23607 31561 sw
rect 2623 28004 15116 28025
rect -15116 27678 -12103 28004
rect -19535 27143 -16883 27678
rect -23307 26434 -21662 27143
tri -21662 26434 -20953 27143 nw
tri -20953 26434 -20244 27143 se
rect -20244 26968 -16883 27143
tri -16883 26968 -16173 27678 nw
tri -16173 26968 -15463 27678 se
rect -15463 27502 -12103 27678
tri -12103 27502 -11601 28004 nw
tri 11601 27502 12103 28004 ne
rect 12103 27502 15116 28004
rect -15463 26968 -12680 27502
rect -20244 26434 -17420 26968
rect -23307 25732 -22364 26434
tri -22364 25732 -21662 26434 nw
tri -21655 25732 -20953 26434 se
rect -20953 26431 -17420 26434
tri -17420 26431 -16883 26968 nw
tri -16710 26431 -16173 26968 se
rect -16173 26925 -12680 26968
tri -12680 26925 -12103 27502 nw
tri -11971 26925 -11394 27502 se
rect -11394 27282 -2268 27502
tri -2268 27282 -2048 27502 sw
rect -11394 26925 -2048 27282
rect -16173 26431 -13174 26925
tri -13174 26431 -12680 26925 nw
tri -12465 26431 -11971 26925 se
rect -11971 26431 -2048 26925
tri -81 26434 987 27502 se
rect 987 26793 11394 27502
tri 11394 26793 12103 27502 sw
tri 12103 26793 12812 27502 ne
rect 12812 27491 15116 27502
tri 15116 27491 15650 28025 sw
tri 15826 27491 16360 28025 ne
rect 16360 27491 19362 28025
rect 12812 26793 15650 27491
rect 987 26434 12103 26793
rect -20953 25732 -18119 26431
tri -18119 25732 -17420 26431 nw
tri -17409 25732 -16710 26431 se
rect -16710 25732 -13873 26431
tri -13873 25732 -13174 26431 nw
tri -13164 25732 -12465 26431 se
rect -12465 25732 -2048 26431
rect -23307 25323 -23073 25732
tri -29436 22196 -26309 25323 se
rect -26309 25023 -23073 25323
tri -23073 25023 -22364 25732 nw
tri -22364 25023 -21655 25732 se
rect -21655 25023 -18829 25732
rect -26309 24316 -23780 25023
tri -23780 24316 -23073 25023 nw
tri -23071 24316 -22364 25023 se
rect -22364 25022 -18829 25023
tri -18829 25022 -18119 25732 nw
tri -18119 25022 -17409 25732 se
rect -17409 25023 -14582 25732
tri -14582 25023 -13873 25732 nw
tri -13873 25023 -13164 25732 se
rect -13164 25222 -2048 25732
rect -13164 25023 -2268 25222
rect -17409 25022 -15116 25023
rect -22364 24489 -19362 25022
tri -19362 24489 -18829 25022 nw
tri -18652 24489 -18119 25022 se
rect -18119 24489 -15116 25022
tri -15116 24489 -14582 25023 nw
tri -14407 24489 -13873 25023 se
rect -13873 25002 -2268 25023
tri -2268 25002 -2048 25222 nw
rect -13873 24489 -11066 25002
rect -22364 24316 -19928 24489
rect -26309 23607 -24489 24316
tri -24489 23607 -23780 24316 nw
tri -23780 23607 -23071 24316 se
rect -23071 23923 -19928 24316
tri -19928 23923 -19362 24489 nw
tri -19218 23923 -18652 24489 se
rect -18652 23923 -15682 24489
tri -15682 23923 -15116 24489 nw
tri -14973 23923 -14407 24489 se
rect -14407 24294 -11066 24489
tri -11066 24294 -10358 25002 nw
tri -2015 24500 -81 26434 se
rect -81 26247 12103 26434
tri 12103 26247 12649 26793 sw
tri 12812 26247 13358 26793 ne
rect 13358 26781 15650 26793
tri 15650 26781 16360 27491 sw
tri 16360 26781 17070 27491 ne
rect 17070 27316 19362 27491
tri 19362 27316 20071 28025 sw
tri 20071 27316 20780 28025 ne
rect 20780 27316 23607 28025
rect 17070 26781 20071 27316
rect 13358 26247 16360 26781
rect -81 25538 12649 26247
tri 12649 25538 13358 26247 sw
tri 13358 25538 14067 26247 ne
rect 14067 26071 16360 26247
tri 16360 26071 17070 26781 sw
tri 17070 26071 17780 26781 ne
rect 17780 26607 20071 26781
tri 20071 26607 20780 27316 sw
tri 20780 26607 21489 27316 ne
rect 21489 26607 23607 27316
rect 17780 26071 20780 26607
rect 14067 25732 17070 26071
tri 17070 25732 17409 26071 sw
tri 17780 25732 18119 26071 ne
rect 18119 25900 20780 26071
tri 20780 25900 21487 26607 sw
tri 21489 25900 22196 26607 ne
rect 22196 25900 23607 26607
rect 18119 25732 21487 25900
rect 14067 25538 17409 25732
rect -81 25002 13358 25538
tri -10356 24294 -10150 24500 se
rect -10150 24294 -81 24500
rect -14407 23923 -11675 24294
rect -23071 23607 -20606 23923
rect -26309 22898 -25198 23607
tri -25198 22898 -24489 23607 nw
tri -24489 22898 -23780 23607 se
rect -23780 23245 -20606 23607
tri -20606 23245 -19928 23923 nw
tri -19896 23245 -19218 23923 se
rect -19218 23245 -16360 23923
tri -16360 23245 -15682 23923 nw
tri -15651 23245 -14973 23923 se
rect -14973 23685 -11675 23923
tri -11675 23685 -11066 24294 nw
tri -10965 23685 -10356 24294 se
rect -10356 23685 -81 24294
rect -14973 23245 -12289 23685
rect -23780 22898 -21274 23245
rect -26309 22196 -25900 22898
tri -25900 22196 -25198 22898 nw
tri -25191 22196 -24489 22898 se
rect -24489 22577 -21274 22898
tri -21274 22577 -20606 23245 nw
tri -20564 22577 -19896 23245 se
rect -19896 22577 -17028 23245
tri -17028 22577 -16360 23245 nw
tri -16319 22577 -15651 23245 se
rect -15651 23071 -12289 23245
tri -12289 23071 -11675 23685 nw
tri -11579 23071 -10965 23685 se
rect -10965 23071 -81 23685
rect -15651 22577 -12996 23071
rect -24489 22196 -21655 22577
tri -21655 22196 -21274 22577 nw
tri -20945 22196 -20564 22577 se
rect -20564 22196 -17603 22577
tri -32972 18660 -29436 22196 se
rect -29436 21487 -26609 22196
tri -26609 21487 -25900 22196 nw
tri -25900 21487 -25191 22196 se
rect -25191 21487 -22365 22196
rect -29436 20780 -27316 21487
tri -27316 20780 -26609 21487 nw
tri -26607 20780 -25900 21487 se
rect -25900 21486 -22365 21487
tri -22365 21486 -21655 22196 nw
tri -21655 21486 -20945 22196 se
rect -20945 22002 -17603 22196
tri -17603 22002 -17028 22577 nw
tri -16894 22002 -16319 22577 se
rect -16319 22364 -12996 22577
tri -12996 22364 -12289 23071 nw
tri -12286 22364 -11579 23071 se
rect -11579 22898 -81 23071
tri -81 22898 2023 25002 nw
tri 10358 24500 10860 25002 ne
rect 10860 24829 13358 25002
tri 13358 24829 14067 25538 sw
tri 14067 24829 14776 25538 ne
rect 14776 25022 17409 25538
tri 17409 25022 18119 25732 sw
tri 18119 25022 18829 25732 ne
rect 18829 25198 21487 25732
tri 21487 25198 22189 25900 sw
tri 22196 25198 22898 25900 ne
rect 22898 25198 23607 25900
rect 18829 25022 22189 25198
rect 14776 24829 18119 25022
rect 10860 24500 14067 24829
tri 2403 24280 2623 24500 se
rect 2623 24280 10150 24500
rect 2403 23966 10150 24280
tri 10150 23966 10684 24500 sw
tri 10860 23966 11394 24500 ne
rect 11394 24489 14067 24500
tri 14067 24489 14407 24829 sw
tri 14776 24489 15116 24829 ne
rect 15116 24489 18119 24829
tri 18119 24489 18652 25022 sw
tri 18829 24489 19362 25022 ne
rect 19362 24489 22189 25022
tri 22189 24489 22898 25198 sw
tri 22898 24489 23607 25198 ne
tri 23607 24489 27143 28025 sw
rect 11394 23966 14407 24489
rect 2403 23432 10684 23966
tri 10684 23432 11218 23966 sw
tri 11394 23432 11928 23966 ne
rect 11928 23780 14407 23966
tri 14407 23780 15116 24489 sw
tri 15116 23780 15825 24489 ne
rect 15825 23955 18652 24489
tri 18652 23955 19186 24489 sw
tri 19362 23955 19896 24489 ne
rect 19896 23955 22898 24489
rect 15825 23780 19186 23955
rect 11928 23432 15116 23780
rect 2403 22898 11218 23432
tri 11218 22898 11752 23432 sw
tri 11928 22898 12462 23432 ne
rect 12462 23245 15116 23432
tri 15116 23245 15651 23780 sw
tri 15825 23245 16360 23780 ne
rect 16360 23245 19186 23780
tri 19186 23245 19896 23955 sw
tri 19896 23245 20606 23955 ne
rect 20606 23780 22898 23955
tri 22898 23780 23607 24489 sw
tri 23607 23780 24316 24489 ne
rect 24316 23780 27143 24489
rect 20606 23245 23607 23780
rect 12462 22898 15651 23245
rect -11579 22364 -979 22898
rect -16319 22002 -13686 22364
rect -20945 21487 -18118 22002
tri -18118 21487 -17603 22002 nw
tri -17409 21487 -16894 22002 se
rect -16894 21674 -13686 22002
tri -13686 21674 -12996 22364 nw
tri -12648 22002 -12286 22364 se
rect -12286 22002 -979 22364
tri -12976 21674 -12648 22002 se
rect -12648 22000 -979 22002
tri -979 22000 -81 22898 nw
rect 2403 22220 11752 22898
tri 2403 22000 2623 22220 ne
rect 2623 22196 11752 22220
tri 11752 22196 12454 22898 sw
tri 12462 22196 13164 22898 ne
rect 13164 22711 15651 22898
tri 15651 22711 16185 23245 sw
tri 16360 22711 16894 23245 ne
rect 16894 22711 19896 23245
rect 13164 22196 16185 22711
rect 2623 22002 12454 22196
tri 12454 22002 12648 22196 sw
tri 13164 22002 13358 22196 ne
rect 13358 22002 16185 22196
tri 16185 22002 16894 22711 sw
tri 16894 22002 17603 22711 ne
rect 17603 22535 19896 22711
tri 19896 22535 20606 23245 sw
tri 20606 22535 21316 23245 ne
rect 21316 23071 23607 23245
tri 23607 23071 24316 23780 sw
tri 24316 23071 25025 23780 ne
rect 25025 23071 27143 23780
rect 21316 22535 24316 23071
rect 17603 22196 20606 22535
tri 20606 22196 20945 22535 sw
tri 21316 22196 21655 22535 ne
rect 21655 22364 24316 22535
tri 24316 22364 25023 23071 sw
tri 25025 22364 25732 23071 ne
rect 25732 22364 27143 23071
rect 21655 22196 25023 22364
rect 17603 22002 20945 22196
rect 2623 22000 12648 22002
rect -16894 21487 -14396 21674
rect -20945 21486 -18652 21487
rect -25900 20953 -22898 21486
tri -22898 20953 -22365 21486 nw
tri -22188 20953 -21655 21486 se
rect -21655 20953 -18652 21486
tri -18652 20953 -18118 21487 nw
tri -17943 20953 -17409 21487 se
rect -17409 20964 -14396 21487
tri -14396 20964 -13686 21674 nw
tri -13686 20964 -12976 21674 se
rect -12976 20964 -12648 21674
rect -17409 20953 -14930 20964
rect -25900 20780 -23245 20953
rect -29436 20071 -28025 20780
tri -28025 20071 -27316 20780 nw
tri -27316 20071 -26607 20780 se
rect -26607 20606 -23245 20780
tri -23245 20606 -22898 20953 nw
tri -22535 20606 -22188 20953 se
rect -22188 20606 -19175 20953
rect -26607 20071 -23955 20606
rect -29436 19362 -28734 20071
tri -28734 19362 -28025 20071 nw
tri -28025 19362 -27316 20071 se
rect -27316 19896 -23955 20071
tri -23955 19896 -23245 20606 nw
tri -23245 19896 -22535 20606 se
rect -22535 20430 -19175 20606
tri -19175 20430 -18652 20953 nw
tri -18466 20430 -17943 20953 se
rect -17943 20430 -14930 20953
tri -14930 20430 -14396 20964 nw
tri -14220 20430 -13686 20964 se
rect -13686 20430 -12648 20964
rect -22535 19896 -19709 20430
tri -19709 19896 -19175 20430 nw
tri -19000 19896 -18466 20430 se
rect -18466 19896 -15464 20430
tri -15464 19896 -14930 20430 nw
tri -14754 19896 -14220 20430 se
rect -14220 19896 -12648 20430
rect -27316 19362 -24489 19896
tri -24489 19362 -23955 19896 nw
tri -23779 19362 -23245 19896 se
rect -23245 19362 -20243 19896
tri -20243 19362 -19709 19896 nw
tri -19534 19362 -19000 19896 se
rect -19000 19362 -15998 19896
tri -15998 19362 -15464 19896 nw
tri -15288 19362 -14754 19896 se
rect -14754 19362 -12648 19896
tri -29436 18660 -28734 19362 nw
tri -28727 18660 -28025 19362 se
rect -28025 18660 -25191 19362
tri -25191 18660 -24489 19362 nw
tri -24481 18660 -23779 19362 se
rect -23779 18660 -20945 19362
tri -20945 18660 -20243 19362 nw
tri -20236 18660 -19534 19362 se
rect -19534 18660 -16700 19362
tri -16700 18660 -15998 19362 nw
tri -15990 18660 -15288 19362 se
rect -15288 18660 -12648 19362
tri -36508 15124 -32972 18660 se
rect -32972 17951 -30145 18660
tri -30145 17951 -29436 18660 nw
tri -29436 17951 -28727 18660 se
rect -28727 17951 -25901 18660
rect -32972 17244 -30852 17951
tri -30852 17244 -30145 17951 nw
tri -30143 17244 -29436 17951 se
rect -29436 17950 -25901 17951
tri -25901 17950 -25191 18660 nw
tri -25191 17950 -24481 18660 se
rect -24481 17951 -21654 18660
tri -21654 17951 -20945 18660 nw
tri -20945 17951 -20236 18660 se
rect -20236 18138 -17222 18660
tri -17222 18138 -16700 18660 nw
tri -16512 18138 -15990 18660 se
rect -15990 18466 -12648 18660
tri -12648 18466 -9114 22000 nw
tri 9114 18466 12648 22000 ne
tri 12648 21468 13182 22002 sw
tri 13358 21468 13892 22002 ne
rect 13892 21468 16894 22002
rect 12648 20758 13182 21468
tri 13182 20758 13892 21468 sw
tri 13892 20758 14602 21468 ne
rect 14602 21293 16894 21468
tri 16894 21293 17603 22002 sw
tri 17603 21293 18312 22002 ne
rect 18312 21486 20945 22002
tri 20945 21486 21655 22196 sw
tri 21655 21486 22365 22196 ne
rect 22365 21662 25023 22196
tri 25023 21662 25725 22364 sw
tri 25732 21662 26434 22364 ne
rect 26434 21662 27143 22364
rect 22365 21486 25725 21662
rect 18312 21293 21655 21486
rect 14602 20953 17603 21293
tri 17603 20953 17943 21293 sw
tri 18312 20953 18652 21293 ne
rect 18652 20953 21655 21293
tri 21655 20953 22188 21486 sw
tri 22365 20953 22898 21486 ne
rect 22898 20953 25725 21486
tri 25725 20953 26434 21662 sw
tri 26434 20953 27143 21662 ne
tri 27143 20953 30679 24489 sw
rect 14602 20758 17943 20953
rect 12648 20048 13892 20758
tri 13892 20048 14602 20758 sw
tri 14602 20048 15312 20758 ne
rect 15312 20244 17943 20758
tri 17943 20244 18652 20953 sw
tri 18652 20244 19361 20953 ne
rect 19361 20419 22188 20953
tri 22188 20419 22722 20953 sw
tri 22898 20419 23432 20953 ne
rect 23432 20419 26434 20953
rect 19361 20244 22722 20419
rect 15312 20048 18652 20244
rect 12648 19362 14602 20048
tri 14602 19362 15288 20048 sw
tri 15312 19362 15998 20048 ne
rect 15998 19709 18652 20048
tri 18652 19709 19187 20244 sw
tri 19361 19709 19896 20244 ne
rect 19896 19709 22722 20244
tri 22722 19709 23432 20419 sw
tri 23432 19709 24142 20419 ne
rect 24142 20244 26434 20419
tri 26434 20244 27143 20953 sw
tri 27143 20244 27852 20953 ne
rect 27852 20244 30679 20953
rect 24142 19709 27143 20244
rect 15998 19362 19187 19709
rect 12648 18660 15288 19362
tri 15288 18660 15990 19362 sw
tri 15998 18660 16700 19362 ne
rect 16700 19175 19187 19362
tri 19187 19175 19721 19709 sw
tri 19896 19175 20430 19709 ne
rect 20430 19175 23432 19709
rect 16700 18660 19721 19175
rect 12648 18466 15990 18660
tri 15990 18466 16184 18660 sw
tri 16700 18466 16894 18660 ne
rect 16894 18466 19721 18660
tri 19721 18466 20430 19175 sw
tri 20430 18466 21139 19175 ne
rect 21139 18999 23432 19175
tri 23432 18999 24142 19709 sw
tri 24142 18999 24852 19709 ne
rect 24852 19535 27143 19709
tri 27143 19535 27852 20244 sw
tri 27852 19535 28561 20244 ne
rect 28561 19535 30679 20244
rect 24852 18999 27852 19535
rect 21139 18660 24142 18999
tri 24142 18660 24481 18999 sw
tri 24852 18660 25191 18999 ne
rect 25191 18828 27852 18999
tri 27852 18828 28559 19535 sw
tri 28561 18828 29268 19535 ne
rect 29268 18828 30679 19535
rect 25191 18660 28559 18828
rect 21139 18466 24481 18660
rect -20236 17951 -17932 18138
rect -24481 17950 -22188 17951
rect -29436 17417 -26434 17950
tri -26434 17417 -25901 17950 nw
tri -25724 17417 -25191 17950 se
rect -25191 17417 -22188 17950
tri -22188 17417 -21654 17951 nw
tri -21479 17417 -20945 17951 se
rect -20945 17428 -17932 17951
tri -17932 17428 -17222 18138 nw
tri -17222 17428 -16512 18138 se
rect -16512 17428 -15990 18138
rect -20945 17417 -18466 17428
rect -29436 17244 -26781 17417
rect -32972 16535 -31561 17244
tri -31561 16535 -30852 17244 nw
tri -30852 16535 -30143 17244 se
rect -30143 17070 -26781 17244
tri -26781 17070 -26434 17417 nw
tri -26071 17070 -25724 17417 se
rect -25724 17070 -22711 17417
rect -30143 16535 -27491 17070
rect -32972 15826 -32270 16535
tri -32270 15826 -31561 16535 nw
tri -31561 15826 -30852 16535 se
rect -30852 16360 -27491 16535
tri -27491 16360 -26781 17070 nw
tri -26781 16360 -26071 17070 se
rect -26071 16894 -22711 17070
tri -22711 16894 -22188 17417 nw
tri -22002 16894 -21479 17417 se
rect -21479 16894 -18466 17417
tri -18466 16894 -17932 17428 nw
tri -17756 16894 -17222 17428 se
rect -17222 16894 -15990 17428
rect -26071 16360 -23245 16894
tri -23245 16360 -22711 16894 nw
tri -22536 16360 -22002 16894 se
rect -22002 16360 -19000 16894
tri -19000 16360 -18466 16894 nw
tri -18290 16360 -17756 16894 se
rect -17756 16360 -15990 16894
rect -30852 15826 -28025 16360
tri -28025 15826 -27491 16360 nw
tri -27315 15826 -26781 16360 se
rect -26781 15826 -23779 16360
tri -23779 15826 -23245 16360 nw
tri -23070 15826 -22536 16360 se
rect -22536 15826 -19534 16360
tri -19534 15826 -19000 16360 nw
tri -18824 15826 -18290 16360 se
rect -18290 15826 -15990 16360
tri -32972 15124 -32270 15826 nw
tri -32263 15124 -31561 15826 se
rect -31561 15124 -28727 15826
tri -28727 15124 -28025 15826 nw
tri -28017 15124 -27315 15826 se
rect -27315 15124 -24481 15826
tri -24481 15124 -23779 15826 nw
tri -23772 15124 -23070 15826 se
rect -23070 15124 -20236 15826
tri -20236 15124 -19534 15826 nw
tri -19526 15124 -18824 15826 se
rect -18824 15124 -15990 15826
tri -15990 15124 -12648 18466 nw
rect -36508 14590 -33506 15124
tri -33506 14590 -32972 15124 nw
tri -32797 14590 -32263 15124 se
rect -32263 14590 -29437 15124
rect -36508 -14590 -34008 14590
tri -34008 14088 -33506 14590 nw
tri -33506 13881 -32797 14590 se
rect -32797 14414 -29437 14590
tri -29437 14414 -28727 15124 nw
tri -28727 14414 -28017 15124 se
rect -28017 14415 -25190 15124
tri -25190 14415 -24481 15124 nw
tri -24481 14415 -23772 15124 se
rect -23772 14602 -20758 15124
tri -20758 14602 -20236 15124 nw
tri -20048 14602 -19526 15124 se
rect -19526 14602 -19513 15124
rect -23772 14415 -21468 14602
rect -28017 14414 -25724 14415
rect -32797 13881 -29970 14414
tri -29970 13881 -29437 14414 nw
tri -29260 13881 -28727 14414 se
rect -28727 13881 -25724 14414
tri -25724 13881 -25190 14415 nw
tri -25015 13881 -24481 14415 se
rect -24481 13892 -21468 14415
tri -21468 13892 -20758 14602 nw
tri -20758 13892 -20048 14602 se
rect -20048 13892 -19513 14602
rect -24481 13881 -22002 13892
rect -33506 13534 -30317 13881
tri -30317 13534 -29970 13881 nw
tri -29607 13534 -29260 13881 se
rect -29260 13534 -26247 13881
rect -33506 -13347 -31006 13534
tri -31006 12845 -30317 13534 nw
tri -30296 12845 -29607 13534 se
rect -29607 13358 -26247 13534
tri -26247 13358 -25724 13881 nw
tri -25538 13358 -25015 13881 se
rect -25015 13358 -22002 13881
tri -22002 13358 -21468 13892 nw
tri -21292 13358 -20758 13892 se
rect -20758 13358 -19513 13892
rect -29607 12845 -26781 13358
tri -30504 12637 -30296 12845 se
rect -30296 12824 -26781 12845
tri -26781 12824 -26247 13358 nw
tri -26072 12824 -25538 13358 se
rect -25538 12824 -22536 13358
tri -22536 12824 -22002 13358 nw
tri -21826 12824 -21292 13358 se
rect -21292 12824 -19513 13358
rect -30296 12637 -26968 12824
tri -26968 12637 -26781 12824 nw
tri -26259 12637 -26072 12824 se
rect -26072 12637 -22723 12824
tri -22723 12637 -22536 12824 nw
tri -22013 12637 -21826 12824 se
rect -21826 12637 -19513 12824
rect -30504 12103 -27502 12637
tri -27502 12103 -26968 12637 nw
tri -26793 12103 -26259 12637 se
rect -26259 12103 -23433 12637
rect -30504 -12103 -28004 12103
tri -28004 11601 -27502 12103 nw
tri -27502 11394 -26793 12103 se
rect -26793 11927 -23433 12103
tri -23433 11927 -22723 12637 nw
tri -22723 11927 -22013 12637 se
rect -22013 11927 -19513 12637
rect -26793 11394 -23966 11927
tri -23966 11394 -23433 11927 nw
tri -23256 11394 -22723 11927 se
rect -22723 11601 -19513 11927
tri -19513 11601 -15990 15124 nw
tri 12648 14930 16184 18466 ne
tri 16184 17932 16718 18466 sw
tri 16894 17932 17428 18466 ne
rect 17428 17932 20430 18466
rect 16184 17222 16718 17932
tri 16718 17222 17428 17932 sw
tri 17428 17222 18138 17932 ne
rect 18138 17757 20430 17932
tri 20430 17757 21139 18466 sw
tri 21139 17757 21848 18466 ne
rect 21848 17950 24481 18466
tri 24481 17950 25191 18660 sw
tri 25191 17950 25901 18660 ne
rect 25901 18126 28559 18660
tri 28559 18126 29261 18828 sw
tri 29268 18126 29970 18828 ne
rect 29970 18126 30679 18828
rect 25901 17950 29261 18126
rect 21848 17757 25191 17950
rect 18138 17417 21139 17757
tri 21139 17417 21479 17757 sw
tri 21848 17417 22188 17757 ne
rect 22188 17417 25191 17757
tri 25191 17417 25724 17950 sw
tri 25901 17417 26434 17950 ne
rect 26434 17417 29261 17950
tri 29261 17417 29970 18126 sw
tri 29970 17417 30679 18126 ne
tri 30679 17417 34215 20953 sw
rect 18138 17222 21479 17417
rect 16184 16512 17428 17222
tri 17428 16512 18138 17222 sw
tri 18138 16512 18848 17222 ne
rect 18848 16708 21479 17222
tri 21479 16708 22188 17417 sw
tri 22188 16708 22897 17417 ne
rect 22897 16883 25724 17417
tri 25724 16883 26258 17417 sw
tri 26434 16883 26968 17417 ne
rect 26968 16883 29970 17417
rect 22897 16708 26258 16883
rect 18848 16512 22188 16708
rect 16184 15826 18138 16512
tri 18138 15826 18824 16512 sw
tri 18848 15826 19534 16512 ne
rect 19534 16173 22188 16512
tri 22188 16173 22723 16708 sw
tri 22897 16173 23432 16708 ne
rect 23432 16173 26258 16708
tri 26258 16173 26968 16883 sw
tri 26968 16173 27678 16883 ne
rect 27678 16708 29970 16883
tri 29970 16708 30679 17417 sw
tri 30679 16708 31388 17417 ne
rect 31388 16708 34215 17417
rect 27678 16173 30679 16708
rect 19534 15826 22723 16173
rect 16184 15124 18824 15826
tri 18824 15124 19526 15826 sw
tri 19534 15124 20236 15826 ne
rect 20236 15639 22723 15826
tri 22723 15639 23257 16173 sw
tri 23432 15639 23966 16173 ne
rect 23966 15639 26968 16173
rect 20236 15124 23257 15639
rect 16184 14930 19526 15124
tri 19526 14930 19720 15124 sw
tri 20236 14930 20430 15124 ne
rect 20430 14930 23257 15124
tri 23257 14930 23966 15639 sw
tri 23966 14930 24675 15639 ne
rect 24675 15463 26968 15639
tri 26968 15463 27678 16173 sw
tri 27678 15463 28388 16173 ne
rect 28388 15999 30679 16173
tri 30679 15999 31388 16708 sw
tri 31388 15999 32097 16708 ne
rect 32097 15999 34215 16708
rect 28388 15463 31388 15999
rect 24675 15124 27678 15463
tri 27678 15124 28017 15463 sw
tri 28388 15124 28727 15463 ne
rect 28727 15292 31388 15463
tri 31388 15292 32095 15999 sw
tri 32097 15292 32804 15999 ne
rect 32804 15292 34215 15999
rect 28727 15124 32095 15292
rect 24675 14930 28017 15124
rect -22723 11394 -22000 11601
rect -27502 11066 -24294 11394
tri -24294 11066 -23966 11394 nw
tri -23584 11066 -23256 11394 se
rect -23256 11066 -22000 11394
rect -27502 -10860 -25002 11066
tri -25002 10358 -24294 11066 nw
tri -24292 10358 -23584 11066 se
rect -23584 10358 -22000 11066
tri -24500 10150 -24292 10358 se
rect -24292 10150 -22000 10358
rect -24500 1250 -22000 10150
tri -22000 9114 -19513 11601 nw
tri 16184 11394 19720 14930 ne
tri 19720 14396 20254 14930 sw
tri 20430 14396 20964 14930 ne
rect 20964 14396 23966 14930
rect 19720 13686 20254 14396
tri 20254 13686 20964 14396 sw
tri 20964 13686 21674 14396 ne
rect 21674 14221 23966 14396
tri 23966 14221 24675 14930 sw
tri 24675 14221 25384 14930 ne
rect 25384 14414 28017 14930
tri 28017 14414 28727 15124 sw
tri 28727 14414 29437 15124 ne
rect 29437 14590 32095 15124
tri 32095 14590 32797 15292 sw
tri 32804 14590 33506 15292 ne
rect 33506 15124 34215 15292
tri 34215 15124 36508 17417 sw
rect 33506 14590 36508 15124
rect 29437 14414 32797 14590
rect 25384 14221 28727 14414
rect 21674 13881 24675 14221
tri 24675 13881 25015 14221 sw
tri 25384 13881 25724 14221 ne
rect 25724 13881 28727 14221
tri 28727 13881 29260 14414 sw
tri 29437 13881 29970 14414 ne
rect 29970 13881 32797 14414
tri 32797 13881 33506 14590 sw
tri 33506 14088 34008 14590 ne
rect 21674 13686 25015 13881
rect 19720 12976 20964 13686
tri 20964 12976 21674 13686 sw
tri 21674 12976 22384 13686 ne
rect 22384 13172 25015 13686
tri 25015 13172 25724 13881 sw
tri 25724 13172 26433 13881 ne
rect 26433 13347 29260 13881
tri 29260 13347 29794 13881 sw
tri 29970 13347 30504 13881 ne
rect 30504 13347 33506 13881
rect 26433 13172 29794 13347
rect 22384 12976 25724 13172
rect 19720 12637 21674 12976
tri 21674 12637 22013 12976 sw
tri 22384 12637 22723 12976 ne
rect 22723 12637 25724 12976
tri 25724 12637 26259 13172 sw
tri 26433 12637 26968 13172 ne
rect 26968 12637 29794 13172
tri 29794 12637 30504 13347 sw
tri 30504 12845 31006 13347 ne
rect 19720 11927 22013 12637
tri 22013 11927 22723 12637 sw
tri 22723 11927 23433 12637 ne
rect 23433 12103 26259 12637
tri 26259 12103 26793 12637 sw
tri 26968 12103 27502 12637 ne
rect 27502 12103 30504 12637
rect 23433 11927 26793 12103
rect 19720 11394 22723 11927
tri 22723 11394 23256 11927 sw
tri 23433 11394 23966 11927 ne
rect 23966 11394 26793 11927
tri 26793 11394 27502 12103 sw
tri 27502 11601 28004 12103 ne
tri 19720 9114 22000 11394 ne
rect 22000 10860 23256 11394
tri 23256 10860 23790 11394 sw
tri 23966 10860 24500 11394 ne
rect 24500 10860 27502 11394
rect 22000 10150 23790 10860
tri 23790 10150 24500 10860 sw
tri 24500 10358 25002 10860 ne
rect -24500 -1250 21000 1250
rect -24500 -10150 -22000 -1250
tri -25002 -10860 -24500 -10358 sw
tri -24500 -10860 -23790 -10150 ne
rect -23790 -10860 -22000 -10150
rect -27502 -11394 -24500 -10860
tri -24500 -11394 -23966 -10860 sw
tri -23790 -11394 -23256 -10860 ne
rect -23256 -11394 -22000 -10860
tri -28004 -12103 -27502 -11601 sw
tri -27502 -12103 -26793 -11394 ne
rect -26793 -11927 -23966 -11394
tri -23966 -11927 -23433 -11394 sw
tri -23256 -11927 -22723 -11394 ne
rect -22723 -11927 -22000 -11394
rect -26793 -12103 -23433 -11927
rect -30504 -12637 -27502 -12103
tri -27502 -12637 -26968 -12103 sw
tri -26793 -12637 -26259 -12103 ne
rect -26259 -12637 -23433 -12103
tri -23433 -12637 -22723 -11927 sw
tri -22723 -12637 -22013 -11927 ne
rect -22013 -12637 -22000 -11927
tri -22000 -12637 -18477 -9114 sw
tri 19513 -11601 22000 -9114 se
rect 22000 -10150 24500 10150
rect 22000 -10358 24292 -10150
tri 24292 -10358 24500 -10150 nw
rect 22000 -11066 23584 -10358
tri 23584 -11066 24292 -10358 nw
tri 24294 -11066 25002 -10358 se
rect 25002 -11066 27502 10860
rect 22000 -11601 23049 -11066
tri 23049 -11601 23584 -11066 nw
tri 23759 -11601 24294 -11066 se
rect 24294 -11394 27502 -11066
rect 24294 -11601 26793 -11394
tri -31006 -13347 -30504 -12845 sw
tri -30504 -13347 -29794 -12637 ne
rect -29794 -13172 -26968 -12637
tri -26968 -13172 -26433 -12637 sw
tri -26259 -13172 -25724 -12637 ne
rect -25724 -12845 -22723 -12637
tri -22723 -12845 -22515 -12637 sw
tri -22013 -12845 -21805 -12637 ne
rect -21805 -12845 -18477 -12637
rect -25724 -13172 -22515 -12845
rect -29794 -13347 -26433 -13172
rect -33506 -13881 -30504 -13347
tri -30504 -13881 -29970 -13347 sw
tri -29794 -13881 -29260 -13347 ne
rect -29260 -13881 -26433 -13347
tri -26433 -13881 -25724 -13172 sw
tri -25724 -13881 -25015 -13172 ne
rect -25015 -13358 -22515 -13172
tri -22515 -13358 -22002 -12845 sw
tri -21805 -13358 -21292 -12845 ne
rect -21292 -13358 -18477 -12845
rect -25015 -13881 -22002 -13358
tri -22002 -13881 -21479 -13358 sw
tri -21292 -13881 -20769 -13358 ne
rect -20769 -13881 -18477 -13358
tri -34008 -14590 -33506 -14088 sw
tri -33506 -14590 -32797 -13881 ne
rect -32797 -14414 -29970 -13881
tri -29970 -14414 -29437 -13881 sw
tri -29260 -14414 -28727 -13881 ne
rect -28727 -14221 -25724 -13881
tri -25724 -14221 -25384 -13881 sw
tri -25015 -14221 -24675 -13881 ne
rect -24675 -14221 -21479 -13881
rect -28727 -14414 -25384 -14221
rect -32797 -14590 -29437 -14414
rect -36508 -15124 -33506 -14590
tri -36508 -17417 -34215 -15124 ne
rect -34215 -15292 -33506 -15124
tri -33506 -15292 -32804 -14590 sw
tri -32797 -15292 -32095 -14590 ne
rect -32095 -15124 -29437 -14590
tri -29437 -15124 -28727 -14414 sw
tri -28727 -15124 -28017 -14414 ne
rect -28017 -14930 -25384 -14414
tri -25384 -14930 -24675 -14221 sw
tri -24675 -14930 -23966 -14221 ne
rect -23966 -14396 -21479 -14221
tri -21479 -14396 -20964 -13881 sw
tri -20769 -14396 -20254 -13881 ne
rect -20254 -14396 -18477 -13881
rect -23966 -14930 -20964 -14396
tri -20964 -14930 -20430 -14396 sw
tri -20254 -14930 -19720 -14396 ne
rect -19720 -14930 -18477 -14396
rect -28017 -15124 -24675 -14930
rect -32095 -15292 -28727 -15124
rect -34215 -16001 -32804 -15292
tri -32804 -16001 -32095 -15292 sw
tri -32095 -16001 -31386 -15292 ne
rect -31386 -15826 -28727 -15292
tri -28727 -15826 -28025 -15124 sw
tri -28017 -15826 -27315 -15124 ne
rect -27315 -15639 -24675 -15124
tri -24675 -15639 -23966 -14930 sw
tri -23966 -15639 -23257 -14930 ne
rect -23257 -15292 -20430 -14930
tri -20430 -15292 -20068 -14930 sw
tri -19720 -15292 -19358 -14930 ne
rect -19358 -15292 -18477 -14930
rect -23257 -15639 -20068 -15292
rect -27315 -15826 -23966 -15639
rect -31386 -16001 -28025 -15826
rect -34215 -16708 -32095 -16001
tri -32095 -16708 -31388 -16001 sw
tri -31386 -16708 -30679 -16001 ne
rect -30679 -16173 -28025 -16001
tri -28025 -16173 -27678 -15826 sw
tri -27315 -16173 -26968 -15826 ne
rect -26968 -16173 -23966 -15826
tri -23966 -16173 -23432 -15639 sw
tri -23257 -16173 -22723 -15639 ne
rect -22723 -15826 -20068 -15639
tri -20068 -15826 -19534 -15292 sw
tri -19358 -15826 -18824 -15292 ne
rect -18824 -15826 -18477 -15292
rect -22723 -16173 -19534 -15826
rect -30679 -16708 -27678 -16173
rect -34215 -17417 -31388 -16708
tri -31388 -17417 -30679 -16708 sw
tri -30679 -17417 -29970 -16708 ne
rect -29970 -16883 -27678 -16708
tri -27678 -16883 -26968 -16173 sw
tri -26968 -16883 -26258 -16173 ne
rect -26258 -16708 -23432 -16173
tri -23432 -16708 -22897 -16173 sw
tri -22723 -16708 -22188 -16173 ne
rect -22188 -16360 -19534 -16173
tri -19534 -16360 -19000 -15826 sw
tri -18824 -16173 -18477 -15826 ne
tri -18477 -16173 -14941 -12637 sw
tri 17026 -14088 19513 -11601 se
rect 19513 -11927 22723 -11601
tri 22723 -11927 23049 -11601 nw
tri 23433 -11927 23759 -11601 se
rect 23759 -11927 26793 -11601
rect 19513 -12637 22013 -11927
tri 22013 -12637 22723 -11927 nw
tri 22723 -12637 23433 -11927 se
rect 23433 -12103 26793 -11927
tri 26793 -12103 27502 -11394 nw
tri 27502 -12103 28004 -11601 se
rect 28004 -12103 30504 12103
rect 23433 -12637 26259 -12103
tri 26259 -12637 26793 -12103 nw
tri 26968 -12637 27502 -12103 se
rect 27502 -12637 30504 -12103
rect 19513 -12845 21805 -12637
tri 21805 -12845 22013 -12637 nw
tri 22515 -12845 22723 -12637 se
rect 22723 -12845 26051 -12637
tri 26051 -12845 26259 -12637 nw
tri 26760 -12845 26968 -12637 se
rect 26968 -12845 30296 -12637
tri 30296 -12845 30504 -12637 nw
rect 19513 -13358 21292 -12845
tri 21292 -13358 21805 -12845 nw
tri 22002 -13358 22515 -12845 se
rect 22515 -13358 25538 -12845
tri 25538 -13358 26051 -12845 nw
tri 26247 -13358 26760 -12845 se
rect 26760 -13358 29607 -12845
rect 19513 -13892 20758 -13358
tri 20758 -13892 21292 -13358 nw
tri 21468 -13892 22002 -13358 se
rect 22002 -13892 24829 -13358
rect 19513 -14088 20048 -13892
tri -18477 -16360 -18290 -16173 ne
rect -18290 -16360 -14941 -16173
rect -22188 -16708 -19000 -16360
rect -26258 -16883 -22897 -16708
rect -29970 -17417 -26968 -16883
tri -26968 -17417 -26434 -16883 sw
tri -26258 -17417 -25724 -16883 ne
rect -25724 -17417 -22897 -16883
tri -22897 -17417 -22188 -16708 sw
tri -22188 -17417 -21479 -16708 ne
rect -21479 -16894 -19000 -16708
tri -19000 -16894 -18466 -16360 sw
tri -18290 -16894 -17756 -16360 ne
rect -17756 -16894 -14941 -16360
rect -21479 -17417 -18466 -16894
tri -18466 -17417 -17943 -16894 sw
tri -17756 -17417 -17233 -16894 ne
rect -17233 -17417 -14941 -16894
tri -34215 -20953 -30679 -17417 ne
tri -30679 -18126 -29970 -17417 sw
tri -29970 -18126 -29261 -17417 ne
rect -29261 -17950 -26434 -17417
tri -26434 -17950 -25901 -17417 sw
tri -25724 -17950 -25191 -17417 ne
rect -25191 -17757 -22188 -17417
tri -22188 -17757 -21848 -17417 sw
tri -21479 -17757 -21139 -17417 ne
rect -21139 -17757 -17943 -17417
rect -25191 -17950 -21848 -17757
rect -29261 -18126 -25901 -17950
rect -30679 -18828 -29970 -18126
tri -29970 -18828 -29268 -18126 sw
tri -29261 -18828 -28559 -18126 ne
rect -28559 -18660 -25901 -18126
tri -25901 -18660 -25191 -17950 sw
tri -25191 -18660 -24481 -17950 ne
rect -24481 -18466 -21848 -17950
tri -21848 -18466 -21139 -17757 sw
tri -21139 -18466 -20430 -17757 ne
rect -20430 -17932 -17943 -17757
tri -17943 -17932 -17428 -17417 sw
tri -17233 -17932 -16718 -17417 ne
rect -16718 -17932 -14941 -17417
rect -20430 -18466 -17428 -17932
tri -17428 -18466 -16894 -17932 sw
tri -16718 -18466 -16184 -17932 ne
rect -16184 -18466 -14941 -17932
rect -24481 -18660 -21139 -18466
rect -28559 -18828 -25191 -18660
rect -30679 -19537 -29268 -18828
tri -29268 -19537 -28559 -18828 sw
tri -28559 -19537 -27850 -18828 ne
rect -27850 -19362 -25191 -18828
tri -25191 -19362 -24489 -18660 sw
tri -24481 -19362 -23779 -18660 ne
rect -23779 -19175 -21139 -18660
tri -21139 -19175 -20430 -18466 sw
tri -20430 -19175 -19721 -18466 ne
rect -19721 -18828 -16894 -18466
tri -16894 -18828 -16532 -18466 sw
tri -16184 -18828 -15822 -18466 ne
rect -15822 -18828 -14941 -18466
rect -19721 -19175 -16532 -18828
rect -23779 -19362 -20430 -19175
rect -27850 -19537 -24489 -19362
rect -30679 -20244 -28559 -19537
tri -28559 -20244 -27852 -19537 sw
tri -27850 -20244 -27143 -19537 ne
rect -27143 -19709 -24489 -19537
tri -24489 -19709 -24142 -19362 sw
tri -23779 -19709 -23432 -19362 ne
rect -23432 -19709 -20430 -19362
tri -20430 -19709 -19896 -19175 sw
tri -19721 -19709 -19187 -19175 ne
rect -19187 -19362 -16532 -19175
tri -16532 -19362 -15998 -18828 sw
tri -15822 -19362 -15288 -18828 ne
rect -15288 -19362 -14941 -18828
rect -19187 -19709 -15998 -19362
rect -27143 -20244 -24142 -19709
rect -30679 -20953 -27852 -20244
tri -27852 -20953 -27143 -20244 sw
tri -27143 -20953 -26434 -20244 ne
rect -26434 -20419 -24142 -20244
tri -24142 -20419 -23432 -19709 sw
tri -23432 -20419 -22722 -19709 ne
rect -22722 -20244 -19896 -19709
tri -19896 -20244 -19361 -19709 sw
tri -19187 -20244 -18652 -19709 ne
rect -18652 -19896 -15998 -19709
tri -15998 -19896 -15464 -19362 sw
tri -15288 -19709 -14941 -19362 ne
tri -14941 -19709 -11405 -16173 sw
tri 13686 -17428 17026 -14088 se
rect 17026 -14602 20048 -14088
tri 20048 -14602 20758 -13892 nw
tri 20758 -14602 21468 -13892 se
rect 21468 -14067 24829 -13892
tri 24829 -14067 25538 -13358 nw
tri 25538 -14067 26247 -13358 se
rect 26247 -13534 29607 -13358
tri 29607 -13534 30296 -12845 nw
tri 30317 -13534 31006 -12845 se
rect 31006 -13534 33506 13347
rect 34008 5500 36508 14590
rect 34008 3000 37508 5500
rect 26247 -14067 29053 -13534
rect 21468 -14415 24481 -14067
tri 24481 -14415 24829 -14067 nw
tri 25190 -14415 25538 -14067 se
rect 25538 -14088 29053 -14067
tri 29053 -14088 29607 -13534 nw
tri 29763 -14088 30317 -13534 se
rect 30317 -13881 33506 -13534
rect 30317 -14088 32797 -13881
rect 25538 -14414 28727 -14088
tri 28727 -14414 29053 -14088 nw
tri 29437 -14414 29763 -14088 se
rect 29763 -14414 32797 -14088
rect 25538 -14415 28017 -14414
rect 21468 -14602 23772 -14415
rect 17026 -15292 19358 -14602
tri 19358 -15292 20048 -14602 nw
tri 20068 -15292 20758 -14602 se
rect 20758 -15124 23772 -14602
tri 23772 -15124 24481 -14415 nw
tri 24481 -15124 25190 -14415 se
rect 25190 -15124 28017 -14415
tri 28017 -15124 28727 -14414 nw
tri 28727 -15124 29437 -14414 se
rect 29437 -14590 32797 -14414
tri 32797 -14590 33506 -13881 nw
rect 34008 -5500 37508 -3000
tri 33506 -14590 34008 -14088 se
rect 34008 -14590 36508 -5500
rect 29437 -15124 32095 -14590
rect 20758 -15292 23070 -15124
rect 17026 -15826 18824 -15292
tri 18824 -15826 19358 -15292 nw
tri 19534 -15826 20068 -15292 se
rect 20068 -15826 23070 -15292
tri 23070 -15826 23772 -15124 nw
tri 23779 -15826 24481 -15124 se
rect 24481 -15826 27315 -15124
tri 27315 -15826 28017 -15124 nw
tri 28025 -15826 28727 -15124 se
rect 28727 -15292 32095 -15124
tri 32095 -15292 32797 -14590 nw
tri 32804 -15292 33506 -14590 se
rect 33506 -15124 36508 -14590
rect 33506 -15292 35806 -15124
rect 28727 -15826 31561 -15292
tri 31561 -15826 32095 -15292 nw
tri 32270 -15826 32804 -15292 se
rect 32804 -15826 35806 -15292
tri 35806 -15826 36508 -15124 nw
rect 17026 -16360 18290 -15826
tri 18290 -16360 18824 -15826 nw
tri 19000 -16360 19534 -15826 se
rect 19534 -16360 22536 -15826
tri 22536 -16360 23070 -15826 nw
tri 23245 -16360 23779 -15826 se
rect 23779 -16360 26781 -15826
tri 26781 -16360 27315 -15826 nw
tri 27491 -16360 28025 -15826 se
rect 28025 -16360 30852 -15826
rect 17026 -16894 17756 -16360
tri 17756 -16894 18290 -16360 nw
tri 18466 -16894 19000 -16360 se
rect 19000 -16894 22002 -16360
tri 22002 -16894 22536 -16360 nw
tri 22711 -16894 23245 -16360 se
rect 23245 -16894 26071 -16360
rect 17026 -17428 17222 -16894
tri 17222 -17428 17756 -16894 nw
tri 17932 -17428 18466 -16894 se
rect 18466 -17428 21293 -16894
tri 11405 -19709 13686 -17428 se
rect 13686 -18138 16512 -17428
tri 16512 -18138 17222 -17428 nw
tri 17222 -18138 17932 -17428 se
rect 17932 -17603 21293 -17428
tri 21293 -17603 22002 -16894 nw
tri 22002 -17603 22711 -16894 se
rect 22711 -17070 26071 -16894
tri 26071 -17070 26781 -16360 nw
tri 26781 -17070 27491 -16360 se
rect 27491 -16535 30852 -16360
tri 30852 -16535 31561 -15826 nw
tri 31561 -16535 32270 -15826 se
rect 27491 -17070 30143 -16535
rect 22711 -17603 25361 -17070
rect 17932 -17951 20945 -17603
tri 20945 -17951 21293 -17603 nw
tri 21654 -17951 22002 -17603 se
rect 22002 -17780 25361 -17603
tri 25361 -17780 26071 -17070 nw
tri 26071 -17780 26781 -17070 se
rect 26781 -17244 30143 -17070
tri 30143 -17244 30852 -16535 nw
tri 30852 -17244 31561 -16535 se
rect 31561 -17244 32270 -16535
rect 26781 -17410 29977 -17244
tri 29977 -17410 30143 -17244 nw
tri 30686 -17410 30852 -17244 se
rect 30852 -17410 32270 -17244
rect 26781 -17780 29268 -17410
rect 22002 -17950 25191 -17780
tri 25191 -17950 25361 -17780 nw
tri 25901 -17950 26071 -17780 se
rect 26071 -17950 29268 -17780
rect 22002 -17951 24481 -17950
rect 17932 -18138 20236 -17951
rect 13686 -18828 15822 -18138
tri 15822 -18828 16512 -18138 nw
tri 16532 -18828 17222 -18138 se
rect 17222 -18660 20236 -18138
tri 20236 -18660 20945 -17951 nw
tri 20945 -18660 21654 -17951 se
rect 21654 -18660 24481 -17951
tri 24481 -18660 25191 -17950 nw
tri 25191 -18660 25901 -17950 se
rect 25901 -18119 29268 -17950
tri 29268 -18119 29977 -17410 nw
tri 29977 -18119 30686 -17410 se
rect 30686 -18119 32270 -17410
rect 25901 -18660 28559 -18119
rect 17222 -18828 19534 -18660
rect 13686 -19362 15288 -18828
tri 15288 -19362 15822 -18828 nw
tri 15998 -19362 16532 -18828 se
rect 16532 -19362 19534 -18828
tri 19534 -19362 20236 -18660 nw
tri 20243 -19362 20945 -18660 se
rect 20945 -19362 23779 -18660
tri 23779 -19362 24481 -18660 nw
tri 24489 -19362 25191 -18660 se
rect 25191 -18828 28559 -18660
tri 28559 -18828 29268 -18119 nw
tri 29268 -18828 29977 -18119 se
rect 29977 -18828 32270 -18119
rect 25191 -19362 28025 -18828
tri 28025 -19362 28559 -18828 nw
tri 28734 -19362 29268 -18828 se
rect 29268 -19362 32270 -18828
tri 32270 -19362 35806 -15826 nw
rect 13686 -19709 14754 -19362
tri -14941 -19896 -14754 -19709 ne
rect -14754 -19896 -11405 -19709
rect -18652 -20244 -15464 -19896
rect -22722 -20419 -19361 -20244
rect -26434 -20953 -23432 -20419
tri -23432 -20953 -22898 -20419 sw
tri -22722 -20953 -22188 -20419 ne
rect -22188 -20953 -19361 -20419
tri -19361 -20953 -18652 -20244 sw
tri -18652 -20953 -17943 -20244 ne
rect -17943 -20430 -15464 -20244
tri -15464 -20430 -14930 -19896 sw
tri -14754 -20430 -14220 -19896 ne
rect -14220 -20430 -11405 -19896
rect -17943 -20953 -14930 -20430
tri -14930 -20953 -14407 -20430 sw
tri -14220 -20953 -13697 -20430 ne
rect -13697 -20953 -11405 -20430
tri -30679 -24489 -27143 -20953 ne
tri -27143 -21662 -26434 -20953 sw
tri -26434 -21662 -25725 -20953 ne
rect -25725 -21486 -22898 -20953
tri -22898 -21486 -22365 -20953 sw
tri -22188 -21486 -21655 -20953 ne
rect -21655 -21293 -18652 -20953
tri -18652 -21293 -18312 -20953 sw
tri -17943 -21293 -17603 -20953 ne
rect -17603 -21293 -14407 -20953
rect -21655 -21486 -18312 -21293
rect -25725 -21662 -22365 -21486
rect -27143 -22364 -26434 -21662
tri -26434 -22364 -25732 -21662 sw
tri -25725 -22364 -25023 -21662 ne
rect -25023 -22196 -22365 -21662
tri -22365 -22196 -21655 -21486 sw
tri -21655 -22196 -20945 -21486 ne
rect -20945 -22002 -18312 -21486
tri -18312 -22002 -17603 -21293 sw
tri -17603 -22002 -16894 -21293 ne
rect -16894 -21468 -14407 -21293
tri -14407 -21468 -13892 -20953 sw
tri -13697 -21468 -13182 -20953 ne
rect -13182 -21468 -11405 -20953
rect -16894 -22002 -13892 -21468
tri -13892 -22002 -13358 -21468 sw
tri -13182 -22002 -12648 -21468 ne
rect -12648 -22000 -11405 -21468
tri -11405 -22000 -9114 -19709 sw
tri 9114 -22000 11405 -19709 se
rect 11405 -19896 14754 -19709
tri 14754 -19896 15288 -19362 nw
tri 15464 -19896 15998 -19362 se
rect 15998 -19896 19000 -19362
tri 19000 -19896 19534 -19362 nw
tri 19709 -19896 20243 -19362 se
rect 20243 -19896 23245 -19362
tri 23245 -19896 23779 -19362 nw
tri 23955 -19896 24489 -19362 se
rect 24489 -19896 27316 -19362
rect 11405 -20430 14220 -19896
tri 14220 -20430 14754 -19896 nw
tri 14930 -20430 15464 -19896 se
rect 15464 -20430 18466 -19896
tri 18466 -20430 19000 -19896 nw
tri 19175 -20430 19709 -19896 se
rect 19709 -20430 22535 -19896
rect 11405 -20964 13686 -20430
tri 13686 -20964 14220 -20430 nw
tri 14396 -20964 14930 -20430 se
rect 14930 -20964 17757 -20430
rect 11405 -21674 12976 -20964
tri 12976 -21674 13686 -20964 nw
tri 13686 -21674 14396 -20964 se
rect 14396 -21139 17757 -20964
tri 17757 -21139 18466 -20430 nw
tri 18466 -21139 19175 -20430 se
rect 19175 -20606 22535 -20430
tri 22535 -20606 23245 -19896 nw
tri 23245 -20606 23955 -19896 se
rect 23955 -20071 27316 -19896
tri 27316 -20071 28025 -19362 nw
tri 28025 -20071 28734 -19362 se
rect 23955 -20606 26607 -20071
rect 19175 -21139 21825 -20606
rect 14396 -21487 17409 -21139
tri 17409 -21487 17757 -21139 nw
tri 18118 -21487 18466 -21139 se
rect 18466 -21316 21825 -21139
tri 21825 -21316 22535 -20606 nw
tri 22535 -21316 23245 -20606 se
rect 23245 -20780 26607 -20606
tri 26607 -20780 27316 -20071 nw
tri 27316 -20780 28025 -20071 se
rect 28025 -20780 28734 -20071
rect 23245 -20946 26441 -20780
tri 26441 -20946 26607 -20780 nw
tri 27150 -20946 27316 -20780 se
rect 27316 -20946 28734 -20780
rect 23245 -21316 25732 -20946
rect 18466 -21486 21655 -21316
tri 21655 -21486 21825 -21316 nw
tri 22365 -21486 22535 -21316 se
rect 22535 -21486 25732 -21316
rect 18466 -21487 20945 -21486
rect 14396 -21674 16700 -21487
rect 11405 -22000 12286 -21674
rect -12648 -22002 12286 -22000
rect -20945 -22196 -17603 -22002
rect -25023 -22364 -21655 -22196
rect -27143 -23073 -25732 -22364
tri -25732 -23073 -25023 -22364 sw
tri -25023 -23073 -24314 -22364 ne
rect -24314 -22898 -21655 -22364
tri -21655 -22898 -20953 -22196 sw
tri -20945 -22898 -20243 -22196 ne
rect -20243 -22711 -17603 -22196
tri -17603 -22711 -16894 -22002 sw
tri -16894 -22711 -16185 -22002 ne
rect -16185 -22364 -13358 -22002
tri -13358 -22364 -12996 -22002 sw
tri -12648 -22364 -12286 -22002 ne
rect -12286 -22364 12286 -22002
tri 12286 -22364 12976 -21674 nw
tri 12996 -22364 13686 -21674 se
rect 13686 -22196 16700 -21674
tri 16700 -22196 17409 -21487 nw
tri 17409 -22196 18118 -21487 se
rect 18118 -22196 20945 -21487
tri 20945 -22196 21655 -21486 nw
tri 21655 -22196 22365 -21486 se
rect 22365 -21655 25732 -21486
tri 25732 -21655 26441 -20946 nw
tri 26441 -21655 27150 -20946 se
rect 27150 -21655 28734 -20946
rect 22365 -22196 25023 -21655
rect 13686 -22364 15998 -22196
rect -16185 -22711 -12996 -22364
rect -20243 -22898 -16894 -22711
rect -24314 -23073 -20953 -22898
rect -27143 -23780 -25023 -23073
tri -25023 -23780 -24316 -23073 sw
tri -24314 -23780 -23607 -23073 ne
rect -23607 -23245 -20953 -23073
tri -20953 -23245 -20606 -22898 sw
tri -20243 -23245 -19896 -22898 ne
rect -19896 -23245 -16894 -22898
tri -16894 -23245 -16360 -22711 sw
tri -16185 -23245 -15651 -22711 ne
rect -15651 -22898 -12996 -22711
tri -12996 -22898 -12462 -22364 sw
tri -12286 -22898 -11752 -22364 ne
rect -11752 -22898 11752 -22364
tri 11752 -22898 12286 -22364 nw
tri 12462 -22898 12996 -22364 se
rect 12996 -22898 15998 -22364
tri 15998 -22898 16700 -22196 nw
tri 16707 -22898 17409 -22196 se
rect 17409 -22898 20243 -22196
tri 20243 -22898 20945 -22196 nw
tri 20953 -22898 21655 -22196 se
rect 21655 -22364 25023 -22196
tri 25023 -22364 25732 -21655 nw
tri 25732 -22364 26441 -21655 se
rect 26441 -22364 28734 -21655
rect 21655 -22898 24489 -22364
tri 24489 -22898 25023 -22364 nw
tri 25198 -22898 25732 -22364 se
rect 25732 -22898 28734 -22364
tri 28734 -22898 32270 -19362 nw
rect -15651 -23245 -12462 -22898
rect -23607 -23780 -20606 -23245
rect -27143 -24489 -24316 -23780
tri -24316 -24489 -23607 -23780 sw
tri -23607 -24489 -22898 -23780 ne
rect -22898 -23955 -20606 -23780
tri -20606 -23955 -19896 -23245 sw
tri -19896 -23955 -19186 -23245 ne
rect -19186 -23780 -16360 -23245
tri -16360 -23780 -15825 -23245 sw
tri -15651 -23780 -15116 -23245 ne
rect -15116 -23432 -12462 -23245
tri -12462 -23432 -11928 -22898 sw
tri -11752 -23432 -11218 -22898 ne
rect -11218 -23432 11218 -22898
tri 11218 -23432 11752 -22898 nw
tri 11928 -23432 12462 -22898 se
rect 12462 -23432 15464 -22898
tri 15464 -23432 15998 -22898 nw
tri 16173 -23432 16707 -22898 se
rect 16707 -23432 19709 -22898
tri 19709 -23432 20243 -22898 nw
tri 20419 -23432 20953 -22898 se
rect 20953 -23432 23780 -22898
rect -15116 -23780 -11928 -23432
rect -19186 -23955 -15825 -23780
rect -22898 -24489 -19896 -23955
tri -19896 -24489 -19362 -23955 sw
tri -19186 -24489 -18652 -23955 ne
rect -18652 -24489 -15825 -23955
tri -15825 -24489 -15116 -23780 sw
tri -15116 -24489 -14407 -23780 ne
rect -14407 -23966 -11928 -23780
tri -11928 -23966 -11394 -23432 sw
tri -11218 -23966 -10684 -23432 ne
rect -10684 -23966 10684 -23432
tri 10684 -23966 11218 -23432 nw
tri 11394 -23966 11928 -23432 se
rect 11928 -23966 14930 -23432
tri 14930 -23966 15464 -23432 nw
tri 15639 -23966 16173 -23432 se
rect 16173 -23966 18999 -23432
rect -14407 -24489 -11394 -23966
tri -11394 -24489 -10871 -23966 sw
tri -10684 -24489 -10161 -23966 ne
rect -10161 -24489 10150 -23966
tri -27143 -28025 -23607 -24489 ne
tri -23607 -25198 -22898 -24489 sw
tri -22898 -25198 -22189 -24489 ne
rect -22189 -25022 -19362 -24489
tri -19362 -25022 -18829 -24489 sw
tri -18652 -25022 -18119 -24489 ne
rect -18119 -25002 -15116 -24489
tri -15116 -25002 -14603 -24489 sw
tri -14407 -25002 -13894 -24489 ne
rect -13894 -25002 -10871 -24489
tri -10871 -25002 -10358 -24489 sw
tri -10161 -24500 -10150 -24489 ne
rect -10150 -24500 10150 -24489
tri 10150 -24500 10684 -23966 nw
tri 10860 -24500 11394 -23966 se
rect 11394 -24500 14221 -23966
tri 10358 -25002 10860 -24500 se
rect 10860 -24675 14221 -24500
tri 14221 -24675 14930 -23966 nw
tri 14930 -24675 15639 -23966 se
rect 15639 -24142 18999 -23966
tri 18999 -24142 19709 -23432 nw
tri 19709 -24142 20419 -23432 se
rect 20419 -23607 23780 -23432
tri 23780 -23607 24489 -22898 nw
tri 24489 -23607 25198 -22898 se
rect 20419 -24142 23071 -23607
rect 15639 -24675 18289 -24142
rect 10860 -25002 13873 -24675
rect -18119 -25022 -14603 -25002
rect -22189 -25198 -18829 -25022
rect -23607 -25900 -22898 -25198
tri -22898 -25900 -22196 -25198 sw
tri -22189 -25900 -21487 -25198 ne
rect -21487 -25732 -18829 -25198
tri -18829 -25732 -18119 -25022 sw
tri -18119 -25732 -17409 -25022 ne
rect -17409 -25580 -14603 -25022
tri -14603 -25580 -14025 -25002 sw
tri -13894 -25580 -13316 -25002 ne
rect -13316 -25580 -979 -25002
rect -17409 -25732 -14025 -25580
rect -21487 -25900 -18119 -25732
rect -23607 -26609 -22196 -25900
tri -22196 -26609 -21487 -25900 sw
tri -21487 -26609 -20778 -25900 ne
rect -20778 -26434 -18119 -25900
tri -18119 -26434 -17417 -25732 sw
tri -17409 -26434 -16707 -25732 ne
rect -16707 -26247 -14025 -25732
tri -14025 -26247 -13358 -25580 sw
tri -13316 -26247 -12649 -25580 ne
rect -12649 -26247 -979 -25580
rect -16707 -26434 -13358 -26247
rect -20778 -26609 -17417 -26434
rect -23607 -27316 -21487 -26609
tri -21487 -27316 -20780 -26609 sw
tri -20778 -27316 -20071 -26609 ne
rect -20071 -26926 -17417 -26609
tri -17417 -26926 -16925 -26434 sw
tri -16707 -26926 -16215 -26434 ne
rect -16215 -26926 -13358 -26434
tri -13358 -26926 -12679 -26247 sw
tri -12649 -26926 -11970 -26247 ne
rect -11970 -26926 -979 -26247
rect -20071 -27316 -16925 -26926
rect -23607 -28025 -20780 -27316
tri -20780 -28025 -20071 -27316 sw
tri -20071 -28025 -19362 -27316 ne
rect -19362 -27491 -16925 -27316
tri -16925 -27491 -16360 -26926 sw
tri -16215 -27491 -15650 -26926 ne
rect -15650 -27491 -12679 -26926
rect -19362 -28025 -16360 -27491
tri -16360 -28025 -15826 -27491 sw
tri -15650 -28025 -15116 -27491 ne
rect -15116 -27502 -12679 -27491
tri -12679 -27502 -12103 -26926 sw
tri -11970 -27502 -11394 -26926 ne
rect -11394 -27502 -979 -26926
rect -15116 -28004 -12103 -27502
tri -12103 -28004 -11601 -27502 sw
rect -15116 -28025 -2380 -28004
tri -23607 -31561 -20071 -28025 ne
tri -20071 -28734 -19362 -28025 sw
tri -19362 -28734 -18653 -28025 ne
rect -18653 -28581 -15826 -28025
tri -15826 -28581 -15270 -28025 sw
tri -15116 -28581 -14560 -28025 ne
rect -14560 -28224 -2380 -28025
tri -2380 -28224 -2160 -28004 sw
tri -2015 -28025 -1492 -27502 ne
rect -1492 -28004 -979 -27502
tri -979 -28004 2023 -25002 sw
tri 2291 -25222 2511 -25002 se
rect 2511 -25023 13873 -25002
tri 13873 -25023 14221 -24675 nw
tri 14582 -25023 14930 -24675 se
rect 14930 -24852 18289 -24675
tri 18289 -24852 18999 -24142 nw
tri 18999 -24852 19709 -24142 se
rect 19709 -24316 23071 -24142
tri 23071 -24316 23780 -23607 nw
tri 23780 -24316 24489 -23607 se
rect 24489 -24316 25198 -23607
rect 19709 -24482 22905 -24316
tri 22905 -24482 23071 -24316 nw
tri 23614 -24482 23780 -24316 se
rect 23780 -24482 25198 -24316
rect 19709 -24852 22196 -24482
rect 14930 -25022 18119 -24852
tri 18119 -25022 18289 -24852 nw
tri 18829 -25022 18999 -24852 se
rect 18999 -25022 22196 -24852
rect 14930 -25023 17409 -25022
rect 2511 -25222 13164 -25023
rect 2291 -25732 13164 -25222
tri 13164 -25732 13873 -25023 nw
tri 13873 -25732 14582 -25023 se
rect 14582 -25732 17409 -25023
tri 17409 -25732 18119 -25022 nw
tri 18119 -25732 18829 -25022 se
rect 18829 -25191 22196 -25022
tri 22196 -25191 22905 -24482 nw
tri 22905 -25191 23614 -24482 se
rect 23614 -25191 25198 -24482
rect 18829 -25732 21487 -25191
rect 2291 -26434 12462 -25732
tri 12462 -26434 13164 -25732 nw
tri 13171 -26434 13873 -25732 se
rect 13873 -26434 16707 -25732
tri 16707 -26434 17409 -25732 nw
tri 17417 -26434 18119 -25732 se
rect 18119 -25900 21487 -25732
tri 21487 -25900 22196 -25191 nw
tri 22196 -25900 22905 -25191 se
rect 22905 -25900 25198 -25191
rect 18119 -26434 20953 -25900
tri 20953 -26434 21487 -25900 nw
tri 21662 -26434 22196 -25900 se
rect 22196 -26434 25198 -25900
tri 25198 -26434 28734 -22898 nw
rect 2291 -26968 11928 -26434
tri 11928 -26968 12462 -26434 nw
tri 12637 -26968 13171 -26434 se
rect 13171 -26968 16173 -26434
tri 16173 -26968 16707 -26434 nw
tri 16883 -26968 17417 -26434 se
rect 17417 -26968 20244 -26434
rect 2291 -27282 11394 -26968
tri 2291 -27502 2511 -27282 ne
rect 2511 -27502 11394 -27282
tri 11394 -27502 11928 -26968 nw
tri 12103 -27502 12637 -26968 se
rect 12637 -27502 15463 -26968
tri 11601 -28004 12103 -27502 se
rect 12103 -27678 15463 -27502
tri 15463 -27678 16173 -26968 nw
tri 16173 -27678 16883 -26968 se
rect 16883 -27143 20244 -26968
tri 20244 -27143 20953 -26434 nw
tri 20953 -27143 21662 -26434 se
rect 16883 -27678 19535 -27143
rect 12103 -28004 14753 -27678
rect -1492 -28025 14753 -28004
rect -14560 -28581 -2160 -28224
rect -18653 -28734 -15270 -28581
rect -20071 -29436 -19362 -28734
tri -19362 -29436 -18660 -28734 sw
tri -18653 -29436 -17951 -28734 ne
rect -17951 -29268 -15270 -28734
tri -15270 -29268 -14583 -28581 sw
tri -14560 -29268 -13873 -28581 ne
rect -13873 -29268 -2160 -28581
rect -17951 -29436 -14583 -29268
rect -20071 -30145 -18660 -29436
tri -18660 -30145 -17951 -29436 sw
tri -17951 -30145 -17242 -29436 ne
rect -17242 -29970 -14583 -29436
tri -14583 -29970 -13881 -29268 sw
tri -13873 -29970 -13171 -29268 ne
rect -13171 -29970 -2160 -29268
rect -17242 -30145 -13881 -29970
rect -20071 -30852 -17951 -30145
tri -17951 -30852 -17244 -30145 sw
tri -17242 -30852 -16535 -30145 ne
rect -16535 -30317 -13881 -30145
tri -13881 -30317 -13534 -29970 sw
tri -13171 -30317 -12824 -29970 ne
rect -12824 -30284 -2160 -29970
rect -12824 -30317 -2380 -30284
rect -16535 -30852 -13534 -30317
rect -20071 -31561 -17244 -30852
tri -17244 -31561 -16535 -30852 sw
tri -16535 -31561 -15826 -30852 ne
rect -15826 -31006 -13534 -30852
tri -13534 -31006 -12845 -30317 sw
tri -12824 -30504 -12637 -30317 ne
rect -12637 -30504 -2380 -30317
tri -2380 -30504 -2160 -30284 nw
tri -1492 -30504 987 -28025 ne
rect 987 -28388 14753 -28025
tri 14753 -28388 15463 -27678 nw
tri 15463 -28388 16173 -27678 se
rect 16173 -27852 19535 -27678
tri 19535 -27852 20244 -27143 nw
tri 20244 -27852 20953 -27143 se
rect 20953 -27852 21662 -27143
rect 16173 -28018 19369 -27852
tri 19369 -28018 19535 -27852 nw
tri 20078 -28018 20244 -27852 se
rect 20244 -28018 21662 -27852
rect 16173 -28388 18660 -28018
rect 987 -28558 14583 -28388
tri 14583 -28558 14753 -28388 nw
tri 15293 -28558 15463 -28388 se
rect 15463 -28558 18660 -28388
rect 987 -29268 13873 -28558
tri 13873 -29268 14583 -28558 nw
tri 14583 -29268 15293 -28558 se
rect 15293 -28727 18660 -28558
tri 18660 -28727 19369 -28018 nw
tri 19369 -28727 20078 -28018 se
rect 20078 -28727 21662 -28018
rect 15293 -29268 17951 -28727
rect 987 -29970 13171 -29268
tri 13171 -29970 13873 -29268 nw
tri 13881 -29970 14583 -29268 se
rect 14583 -29436 17951 -29268
tri 17951 -29436 18660 -28727 nw
tri 18660 -29436 19369 -28727 se
rect 19369 -29436 21662 -28727
rect 14583 -29970 17417 -29436
tri 17417 -29970 17951 -29436 nw
tri 18126 -29970 18660 -29436 se
rect 18660 -29970 21662 -29436
tri 21662 -29970 25198 -26434 nw
rect 987 -30504 12637 -29970
tri 12637 -30504 13171 -29970 nw
tri 13347 -30504 13881 -29970 se
rect 13881 -30504 16708 -29970
tri 12845 -31006 13347 -30504 se
rect 13347 -30679 16708 -30504
tri 16708 -30679 17417 -29970 nw
tri 17417 -30679 18126 -29970 se
rect 13347 -31006 15999 -30679
rect -15826 -31561 -979 -31006
tri -20071 -35079 -16553 -31561 ne
rect -16553 -32270 -16535 -31561
tri -16535 -32270 -15826 -31561 sw
tri -15826 -32270 -15117 -31561 ne
rect -15117 -32270 -979 -31561
rect -16553 -32972 -15826 -32270
tri -15826 -32972 -15124 -32270 sw
tri -15117 -32972 -14415 -32270 ne
rect -14415 -32972 -979 -32270
rect -16553 -33506 -15124 -32972
tri -15124 -33506 -14590 -32972 sw
tri -14415 -33506 -13881 -32972 ne
rect -13881 -33506 -979 -32972
rect -16553 -34008 -14590 -33506
tri -14590 -34008 -14088 -33506 sw
tri -2015 -34008 -1513 -33506 ne
rect -1513 -34008 -979 -33506
tri -979 -34008 2023 -31006 sw
tri 2291 -31226 2511 -31006 se
rect 2511 -31226 15999 -31006
rect 2291 -31388 15999 -31226
tri 15999 -31388 16708 -30679 nw
tri 16708 -31388 17417 -30679 se
rect 17417 -31388 18126 -30679
rect 2291 -31554 15833 -31388
tri 15833 -31554 15999 -31388 nw
tri 16542 -31554 16708 -31388 se
rect 16708 -31554 18126 -31388
rect 2291 -32263 15124 -31554
tri 15124 -32263 15833 -31554 nw
tri 15833 -32263 16542 -31554 se
rect 16542 -32263 18126 -31554
rect 2291 -32972 14415 -32263
tri 14415 -32972 15124 -32263 nw
tri 15124 -32972 15833 -32263 se
rect 15833 -32972 18126 -32263
rect 2291 -33286 13881 -32972
tri 2291 -33506 2511 -33286 ne
rect 2511 -33506 13881 -33286
tri 13881 -33506 14415 -32972 nw
tri 14590 -33506 15124 -32972 se
rect 15124 -33506 18126 -32972
tri 18126 -33506 21662 -29970 nw
tri 14088 -34008 14590 -33506 se
rect 14590 -34008 15124 -33506
rect -16553 -34228 -2380 -34008
tri -2380 -34228 -2160 -34008 sw
rect -16553 -35079 -2160 -34228
tri -16553 -36508 -15124 -35079 ne
rect -15124 -36288 -2160 -35079
rect -15124 -36508 -2380 -36288
tri -2380 -36508 -2160 -36288 nw
tri -1513 -36508 987 -34008 ne
rect 987 -36508 15124 -34008
tri 15124 -36508 18126 -33506 nw
<< properties >>
string FIXED_BBOX 0 0 74016 73016
string LEFclass BLOCK
string LEFview TRUE
string gencell sky130_fd_pr__rf_test_coil3
string library sky130
string parameter m=1
string GDS_END 10411016
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10379748
<< end >>
