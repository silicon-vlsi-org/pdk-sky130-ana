magic
tech sky130A
magscale 1 2
timestamp 1746986264
<< nwell >>
rect -10 0 893 1292
<< pmos >>
rect 194 141 224 1151
rect 348 141 378 1151
rect 502 141 532 1151
rect 656 141 686 1151
<< pdiff >>
rect 138 1139 194 1151
rect 138 1105 149 1139
rect 183 1105 194 1139
rect 138 1071 194 1105
rect 138 1037 149 1071
rect 183 1037 194 1071
rect 138 1003 194 1037
rect 138 969 149 1003
rect 183 969 194 1003
rect 138 935 194 969
rect 138 901 149 935
rect 183 901 194 935
rect 138 867 194 901
rect 138 833 149 867
rect 183 833 194 867
rect 138 799 194 833
rect 138 765 149 799
rect 183 765 194 799
rect 138 731 194 765
rect 138 697 149 731
rect 183 697 194 731
rect 138 663 194 697
rect 138 629 149 663
rect 183 629 194 663
rect 138 595 194 629
rect 138 561 149 595
rect 183 561 194 595
rect 138 527 194 561
rect 138 493 149 527
rect 183 493 194 527
rect 138 459 194 493
rect 138 425 149 459
rect 183 425 194 459
rect 138 391 194 425
rect 138 357 149 391
rect 183 357 194 391
rect 138 323 194 357
rect 138 289 149 323
rect 183 289 194 323
rect 138 255 194 289
rect 138 221 149 255
rect 183 221 194 255
rect 138 187 194 221
rect 138 153 149 187
rect 183 153 194 187
rect 138 141 194 153
rect 224 1139 348 1151
rect 224 153 235 1139
rect 337 153 348 1139
rect 224 141 348 153
rect 378 1139 502 1151
rect 378 153 389 1139
rect 491 153 502 1139
rect 378 141 502 153
rect 532 1139 656 1151
rect 532 153 543 1139
rect 645 153 656 1139
rect 532 141 656 153
rect 686 1139 745 1151
rect 686 1105 697 1139
rect 731 1105 745 1139
rect 686 1071 745 1105
rect 686 1037 697 1071
rect 731 1037 745 1071
rect 686 1003 745 1037
rect 686 969 697 1003
rect 731 969 745 1003
rect 686 935 745 969
rect 686 901 697 935
rect 731 901 745 935
rect 686 867 745 901
rect 686 833 697 867
rect 731 833 745 867
rect 686 799 745 833
rect 686 765 697 799
rect 731 765 745 799
rect 686 731 745 765
rect 686 697 697 731
rect 731 697 745 731
rect 686 663 745 697
rect 686 629 697 663
rect 731 629 745 663
rect 686 595 745 629
rect 686 561 697 595
rect 731 561 745 595
rect 686 527 745 561
rect 686 493 697 527
rect 731 493 745 527
rect 686 459 745 493
rect 686 425 697 459
rect 731 425 745 459
rect 686 391 745 425
rect 686 357 697 391
rect 731 357 745 391
rect 686 323 745 357
rect 686 289 697 323
rect 731 289 745 323
rect 686 255 745 289
rect 686 221 697 255
rect 731 221 745 255
rect 686 187 745 221
rect 686 153 697 187
rect 731 153 745 187
rect 686 141 745 153
<< pdiffc >>
rect 149 1105 183 1139
rect 149 1037 183 1071
rect 149 969 183 1003
rect 149 901 183 935
rect 149 833 183 867
rect 149 765 183 799
rect 149 697 183 731
rect 149 629 183 663
rect 149 561 183 595
rect 149 493 183 527
rect 149 425 183 459
rect 149 357 183 391
rect 149 289 183 323
rect 149 221 183 255
rect 149 153 183 187
rect 235 153 337 1139
rect 389 153 491 1139
rect 543 153 645 1139
rect 697 1105 731 1139
rect 697 1037 731 1071
rect 697 969 731 1003
rect 697 901 731 935
rect 697 833 731 867
rect 697 765 731 799
rect 697 697 731 731
rect 697 629 731 663
rect 697 561 731 595
rect 697 493 731 527
rect 697 425 731 459
rect 697 357 731 391
rect 697 289 731 323
rect 697 221 731 255
rect 697 153 731 187
<< nsubdiff >>
rect 26 1105 84 1151
rect 26 1071 38 1105
rect 72 1071 84 1105
rect 26 1037 84 1071
rect 26 1003 38 1037
rect 72 1003 84 1037
rect 26 969 84 1003
rect 26 935 38 969
rect 72 935 84 969
rect 26 901 84 935
rect 26 867 38 901
rect 72 867 84 901
rect 26 833 84 867
rect 26 799 38 833
rect 72 799 84 833
rect 26 765 84 799
rect 26 731 38 765
rect 72 731 84 765
rect 26 697 84 731
rect 26 663 38 697
rect 72 663 84 697
rect 26 629 84 663
rect 26 595 38 629
rect 72 595 84 629
rect 26 561 84 595
rect 26 527 38 561
rect 72 527 84 561
rect 26 493 84 527
rect 26 459 38 493
rect 72 459 84 493
rect 26 425 84 459
rect 26 391 38 425
rect 72 391 84 425
rect 26 357 84 391
rect 26 323 38 357
rect 72 323 84 357
rect 26 289 84 323
rect 26 255 38 289
rect 72 255 84 289
rect 26 221 84 255
rect 26 187 38 221
rect 72 187 84 221
rect 26 141 84 187
rect 799 1105 857 1151
rect 799 1071 811 1105
rect 845 1071 857 1105
rect 799 1037 857 1071
rect 799 1003 811 1037
rect 845 1003 857 1037
rect 799 969 857 1003
rect 799 935 811 969
rect 845 935 857 969
rect 799 901 857 935
rect 799 867 811 901
rect 845 867 857 901
rect 799 833 857 867
rect 799 799 811 833
rect 845 799 857 833
rect 799 765 857 799
rect 799 731 811 765
rect 845 731 857 765
rect 799 697 857 731
rect 799 663 811 697
rect 845 663 857 697
rect 799 629 857 663
rect 799 595 811 629
rect 845 595 857 629
rect 799 561 857 595
rect 799 527 811 561
rect 845 527 857 561
rect 799 493 857 527
rect 799 459 811 493
rect 845 459 857 493
rect 799 425 857 459
rect 799 391 811 425
rect 845 391 857 425
rect 799 357 857 391
rect 799 323 811 357
rect 845 323 857 357
rect 799 289 857 323
rect 799 255 811 289
rect 845 255 857 289
rect 799 221 857 255
rect 799 187 811 221
rect 845 187 857 221
rect 799 141 857 187
<< nsubdiffcont >>
rect 38 1071 72 1105
rect 38 1003 72 1037
rect 38 935 72 969
rect 38 867 72 901
rect 38 799 72 833
rect 38 731 72 765
rect 38 663 72 697
rect 38 595 72 629
rect 38 527 72 561
rect 38 459 72 493
rect 38 391 72 425
rect 38 323 72 357
rect 38 255 72 289
rect 38 187 72 221
rect 811 1071 845 1105
rect 811 1003 845 1037
rect 811 935 845 969
rect 811 867 845 901
rect 811 799 845 833
rect 811 731 845 765
rect 811 663 845 697
rect 811 595 845 629
rect 811 527 845 561
rect 811 459 845 493
rect 811 391 845 425
rect 811 323 845 357
rect 811 255 845 289
rect 811 187 845 221
<< poly >>
rect 194 1246 736 1262
rect 194 1212 210 1246
rect 244 1212 278 1246
rect 312 1212 346 1246
rect 380 1212 414 1246
rect 448 1212 482 1246
rect 516 1212 550 1246
rect 584 1212 618 1246
rect 652 1212 686 1246
rect 720 1212 736 1246
rect 194 1196 736 1212
rect 194 1151 224 1196
rect 348 1151 378 1196
rect 502 1151 532 1196
rect 656 1151 686 1196
rect 194 96 224 141
rect 348 96 378 141
rect 502 96 532 141
rect 656 96 686 141
rect 194 80 736 96
rect 194 46 210 80
rect 244 46 278 80
rect 312 46 346 80
rect 380 46 414 80
rect 448 46 482 80
rect 516 46 550 80
rect 584 46 618 80
rect 652 46 686 80
rect 720 46 736 80
rect 194 30 736 46
<< polycont >>
rect 210 1212 244 1246
rect 278 1212 312 1246
rect 346 1212 380 1246
rect 414 1212 448 1246
rect 482 1212 516 1246
rect 550 1212 584 1246
rect 618 1212 652 1246
rect 686 1212 720 1246
rect 210 46 244 80
rect 278 46 312 80
rect 346 46 380 80
rect 414 46 448 80
rect 482 46 516 80
rect 550 46 584 80
rect 618 46 652 80
rect 686 46 720 80
<< locali >>
rect 244 1212 266 1246
rect 312 1212 338 1246
rect 380 1212 410 1246
rect 448 1212 482 1246
rect 516 1212 550 1246
rect 588 1212 618 1246
rect 660 1212 686 1246
rect 732 1212 736 1246
rect 149 1139 183 1155
rect 38 1059 72 1071
rect 38 987 72 1003
rect 38 915 72 935
rect 38 843 72 867
rect 38 771 72 799
rect 38 699 72 731
rect 38 629 72 663
rect 38 561 72 593
rect 38 493 72 521
rect 38 425 72 449
rect 38 357 72 377
rect 38 289 72 305
rect 38 221 72 233
rect 149 1071 183 1097
rect 149 1003 183 1025
rect 149 935 183 953
rect 149 867 183 881
rect 149 799 183 809
rect 149 731 183 737
rect 149 663 183 665
rect 149 627 183 629
rect 149 555 183 561
rect 149 483 183 493
rect 149 411 183 425
rect 149 339 183 357
rect 149 267 183 289
rect 149 195 183 221
rect 149 137 183 153
rect 233 1139 339 1155
rect 233 1131 235 1139
rect 337 1131 339 1139
rect 233 153 235 161
rect 337 153 339 161
rect 233 137 339 153
rect 387 1139 493 1155
rect 387 1131 389 1139
rect 491 1131 493 1139
rect 387 153 389 161
rect 491 153 493 161
rect 387 137 493 153
rect 541 1139 647 1155
rect 541 1131 543 1139
rect 645 1131 647 1139
rect 541 153 543 161
rect 645 153 647 161
rect 541 137 647 153
rect 697 1139 731 1155
rect 697 1071 731 1097
rect 697 1003 731 1025
rect 697 935 731 953
rect 697 867 731 881
rect 697 799 731 809
rect 697 731 731 737
rect 697 663 731 665
rect 697 627 731 629
rect 697 555 731 561
rect 697 483 731 493
rect 697 411 731 425
rect 697 339 731 357
rect 697 267 731 289
rect 697 195 731 221
rect 811 1059 845 1071
rect 811 987 845 1003
rect 811 915 845 935
rect 811 843 845 867
rect 811 771 845 799
rect 811 699 845 731
rect 811 629 845 663
rect 811 561 845 593
rect 811 493 845 521
rect 811 425 845 449
rect 811 357 845 377
rect 811 289 845 305
rect 811 221 845 233
rect 697 137 731 153
rect 244 46 266 80
rect 312 46 338 80
rect 380 46 410 80
rect 448 46 482 80
rect 516 46 550 80
rect 588 46 618 80
rect 660 46 686 80
rect 732 46 736 80
<< viali >>
rect 194 1212 210 1246
rect 210 1212 228 1246
rect 266 1212 278 1246
rect 278 1212 300 1246
rect 338 1212 346 1246
rect 346 1212 372 1246
rect 410 1212 414 1246
rect 414 1212 444 1246
rect 482 1212 516 1246
rect 554 1212 584 1246
rect 584 1212 588 1246
rect 626 1212 652 1246
rect 652 1212 660 1246
rect 698 1212 720 1246
rect 720 1212 732 1246
rect 38 1105 72 1131
rect 38 1097 72 1105
rect 38 1037 72 1059
rect 38 1025 72 1037
rect 38 969 72 987
rect 38 953 72 969
rect 38 901 72 915
rect 38 881 72 901
rect 38 833 72 843
rect 38 809 72 833
rect 38 765 72 771
rect 38 737 72 765
rect 38 697 72 699
rect 38 665 72 697
rect 38 595 72 627
rect 38 593 72 595
rect 38 527 72 555
rect 38 521 72 527
rect 38 459 72 483
rect 38 449 72 459
rect 38 391 72 411
rect 38 377 72 391
rect 38 323 72 339
rect 38 305 72 323
rect 38 255 72 267
rect 38 233 72 255
rect 38 187 72 195
rect 38 161 72 187
rect 149 1105 183 1131
rect 149 1097 183 1105
rect 149 1037 183 1059
rect 149 1025 183 1037
rect 149 969 183 987
rect 149 953 183 969
rect 149 901 183 915
rect 149 881 183 901
rect 149 833 183 843
rect 149 809 183 833
rect 149 765 183 771
rect 149 737 183 765
rect 149 697 183 699
rect 149 665 183 697
rect 149 595 183 627
rect 149 593 183 595
rect 149 527 183 555
rect 149 521 183 527
rect 149 459 183 483
rect 149 449 183 459
rect 149 391 183 411
rect 149 377 183 391
rect 149 323 183 339
rect 149 305 183 323
rect 149 255 183 267
rect 149 233 183 255
rect 149 187 183 195
rect 149 161 183 187
rect 233 161 235 1131
rect 235 161 337 1131
rect 337 161 339 1131
rect 387 161 389 1131
rect 389 161 491 1131
rect 491 161 493 1131
rect 541 161 543 1131
rect 543 161 645 1131
rect 645 161 647 1131
rect 697 1105 731 1131
rect 697 1097 731 1105
rect 697 1037 731 1059
rect 697 1025 731 1037
rect 697 969 731 987
rect 697 953 731 969
rect 697 901 731 915
rect 697 881 731 901
rect 697 833 731 843
rect 697 809 731 833
rect 697 765 731 771
rect 697 737 731 765
rect 697 697 731 699
rect 697 665 731 697
rect 697 595 731 627
rect 697 593 731 595
rect 697 527 731 555
rect 697 521 731 527
rect 697 459 731 483
rect 697 449 731 459
rect 697 391 731 411
rect 697 377 731 391
rect 697 323 731 339
rect 697 305 731 323
rect 697 255 731 267
rect 697 233 731 255
rect 697 187 731 195
rect 697 161 731 187
rect 811 1105 845 1131
rect 811 1097 845 1105
rect 811 1037 845 1059
rect 811 1025 845 1037
rect 811 969 845 987
rect 811 953 845 969
rect 811 901 845 915
rect 811 881 845 901
rect 811 833 845 843
rect 811 809 845 833
rect 811 765 845 771
rect 811 737 845 765
rect 811 697 845 699
rect 811 665 845 697
rect 811 595 845 627
rect 811 593 845 595
rect 811 527 845 555
rect 811 521 845 527
rect 811 459 845 483
rect 811 449 845 459
rect 811 391 845 411
rect 811 377 845 391
rect 811 323 845 339
rect 811 305 845 323
rect 811 255 845 267
rect 811 233 845 255
rect 811 187 845 195
rect 811 161 845 187
rect 194 46 210 80
rect 210 46 228 80
rect 266 46 278 80
rect 278 46 300 80
rect 338 46 346 80
rect 346 46 372 80
rect 410 46 414 80
rect 414 46 444 80
rect 482 46 516 80
rect 554 46 584 80
rect 584 46 588 80
rect 626 46 652 80
rect 652 46 660 80
rect 698 46 720 80
rect 720 46 732 80
<< metal1 >>
rect 182 1246 744 1258
rect 182 1212 194 1246
rect 228 1212 266 1246
rect 300 1212 338 1246
rect 372 1212 410 1246
rect 444 1212 482 1246
rect 516 1212 554 1246
rect 588 1212 626 1246
rect 660 1212 698 1246
rect 732 1212 744 1246
rect 182 1200 744 1212
rect 140 1148 192 1154
rect 26 1131 84 1143
rect 26 1097 38 1131
rect 72 1097 84 1131
rect 26 1059 84 1097
rect 26 1025 38 1059
rect 72 1025 84 1059
rect 26 987 84 1025
rect 26 953 38 987
rect 72 953 84 987
rect 26 915 84 953
rect 26 881 38 915
rect 72 881 84 915
rect 26 843 84 881
rect 26 809 38 843
rect 72 809 84 843
rect 26 771 84 809
rect 26 737 38 771
rect 72 737 84 771
rect 26 699 84 737
rect 26 665 38 699
rect 72 665 84 699
rect 26 627 84 665
rect 26 593 38 627
rect 72 593 84 627
rect 26 555 84 593
rect 26 521 38 555
rect 72 521 84 555
rect 26 483 84 521
rect 26 449 38 483
rect 72 449 84 483
rect 26 411 84 449
rect 26 377 38 411
rect 72 377 84 411
rect 26 339 84 377
rect 26 305 38 339
rect 72 305 84 339
rect 26 267 84 305
rect 26 233 38 267
rect 72 233 84 267
rect 26 195 84 233
rect 26 161 38 195
rect 72 161 84 195
rect 26 149 84 161
rect 382 1149 498 1155
rect 192 1096 195 1143
rect 140 1084 195 1096
rect 192 1032 195 1084
rect 140 1025 149 1032
rect 183 1025 195 1032
rect 140 1020 195 1025
rect 192 968 195 1020
rect 140 956 149 968
rect 183 956 195 968
rect 192 904 195 956
rect 140 881 149 904
rect 183 881 195 904
rect 140 843 195 881
rect 140 809 149 843
rect 183 809 195 843
rect 140 771 195 809
rect 140 737 149 771
rect 183 737 195 771
rect 140 699 195 737
rect 140 665 149 699
rect 183 665 195 699
rect 140 627 195 665
rect 140 593 149 627
rect 183 593 195 627
rect 140 555 195 593
rect 140 521 149 555
rect 183 521 195 555
rect 140 483 195 521
rect 140 449 149 483
rect 183 449 195 483
rect 140 411 195 449
rect 140 388 149 411
rect 183 388 195 411
rect 192 336 195 388
rect 140 324 149 336
rect 183 324 195 336
rect 192 272 195 324
rect 140 267 195 272
rect 140 260 149 267
rect 183 260 195 267
rect 192 208 195 260
rect 140 196 195 208
rect 192 149 195 196
rect 223 1131 349 1143
rect 223 864 233 1131
rect 339 864 349 1131
rect 223 428 228 864
rect 344 428 349 864
rect 223 161 233 428
rect 339 161 349 428
rect 223 149 349 161
rect 377 905 382 1143
rect 688 1149 740 1155
rect 498 905 503 1143
rect 377 161 387 905
rect 493 161 503 905
rect 377 149 503 161
rect 531 1131 657 1143
rect 531 864 541 1131
rect 647 864 657 1131
rect 531 428 536 864
rect 652 428 657 864
rect 531 161 541 428
rect 647 161 657 428
rect 531 149 657 161
rect 685 1097 688 1143
rect 740 1097 743 1143
rect 685 1085 743 1097
rect 685 1033 688 1085
rect 740 1033 743 1085
rect 685 1025 697 1033
rect 731 1025 743 1033
rect 685 1021 743 1025
rect 685 969 688 1021
rect 740 969 743 1021
rect 685 957 697 969
rect 731 957 743 969
rect 685 905 688 957
rect 740 905 743 957
rect 685 881 697 905
rect 731 881 743 905
rect 685 843 743 881
rect 685 809 697 843
rect 731 809 743 843
rect 685 771 743 809
rect 685 737 697 771
rect 731 737 743 771
rect 685 699 743 737
rect 685 665 697 699
rect 731 665 743 699
rect 685 627 743 665
rect 685 593 697 627
rect 731 593 743 627
rect 685 555 743 593
rect 685 521 697 555
rect 731 521 743 555
rect 685 483 743 521
rect 685 449 697 483
rect 731 449 743 483
rect 685 411 743 449
rect 685 388 697 411
rect 731 388 743 411
rect 685 336 688 388
rect 740 336 743 388
rect 685 324 697 336
rect 731 324 743 336
rect 685 272 688 324
rect 740 272 743 324
rect 685 267 743 272
rect 685 260 697 267
rect 731 260 743 267
rect 685 208 688 260
rect 740 208 743 260
rect 685 196 743 208
rect 685 149 688 196
rect 140 138 192 144
rect 740 149 743 196
rect 799 1131 857 1143
rect 799 1097 811 1131
rect 845 1097 857 1131
rect 799 1059 857 1097
rect 799 1025 811 1059
rect 845 1025 857 1059
rect 799 987 857 1025
rect 799 953 811 987
rect 845 953 857 987
rect 799 915 857 953
rect 799 881 811 915
rect 845 881 857 915
rect 799 843 857 881
rect 799 809 811 843
rect 845 809 857 843
rect 799 771 857 809
rect 799 737 811 771
rect 845 737 857 771
rect 799 699 857 737
rect 799 665 811 699
rect 845 665 857 699
rect 799 627 857 665
rect 799 593 811 627
rect 845 593 857 627
rect 799 555 857 593
rect 799 521 811 555
rect 845 521 857 555
rect 799 483 857 521
rect 799 449 811 483
rect 845 449 857 483
rect 799 411 857 449
rect 799 377 811 411
rect 845 377 857 411
rect 799 339 857 377
rect 799 305 811 339
rect 845 305 857 339
rect 799 267 857 305
rect 799 233 811 267
rect 845 233 857 267
rect 799 195 857 233
rect 799 161 811 195
rect 845 161 857 195
rect 799 149 857 161
rect 688 138 740 144
rect 182 80 744 92
rect 182 46 194 80
rect 228 46 266 80
rect 300 46 338 80
rect 372 46 410 80
rect 444 46 482 80
rect 516 46 554 80
rect 588 46 626 80
rect 660 46 698 80
rect 732 46 744 80
rect 182 34 744 46
<< via1 >>
rect 140 1131 192 1148
rect 140 1097 149 1131
rect 149 1097 183 1131
rect 183 1097 192 1131
rect 140 1096 192 1097
rect 140 1059 192 1084
rect 140 1032 149 1059
rect 149 1032 183 1059
rect 183 1032 192 1059
rect 140 987 192 1020
rect 140 968 149 987
rect 149 968 183 987
rect 183 968 192 987
rect 140 953 149 956
rect 149 953 183 956
rect 183 953 192 956
rect 140 915 192 953
rect 140 904 149 915
rect 149 904 183 915
rect 183 904 192 915
rect 140 377 149 388
rect 149 377 183 388
rect 183 377 192 388
rect 140 339 192 377
rect 140 336 149 339
rect 149 336 183 339
rect 183 336 192 339
rect 140 305 149 324
rect 149 305 183 324
rect 183 305 192 324
rect 140 272 192 305
rect 140 233 149 260
rect 149 233 183 260
rect 183 233 192 260
rect 140 208 192 233
rect 140 195 192 196
rect 140 161 149 195
rect 149 161 183 195
rect 183 161 192 195
rect 140 144 192 161
rect 228 428 233 864
rect 233 428 339 864
rect 339 428 344 864
rect 382 1131 498 1149
rect 382 905 387 1131
rect 387 905 493 1131
rect 493 905 498 1131
rect 536 428 541 864
rect 541 428 647 864
rect 647 428 652 864
rect 688 1131 740 1149
rect 688 1097 697 1131
rect 697 1097 731 1131
rect 731 1097 740 1131
rect 688 1059 740 1085
rect 688 1033 697 1059
rect 697 1033 731 1059
rect 731 1033 740 1059
rect 688 987 740 1021
rect 688 969 697 987
rect 697 969 731 987
rect 731 969 740 987
rect 688 953 697 957
rect 697 953 731 957
rect 731 953 740 957
rect 688 915 740 953
rect 688 905 697 915
rect 697 905 731 915
rect 731 905 740 915
rect 688 377 697 388
rect 697 377 731 388
rect 731 377 740 388
rect 688 339 740 377
rect 688 336 697 339
rect 697 336 731 339
rect 731 336 740 339
rect 688 305 697 324
rect 697 305 731 324
rect 731 305 740 324
rect 688 272 740 305
rect 688 233 697 260
rect 697 233 731 260
rect 731 233 740 260
rect 688 208 740 233
rect 688 195 740 196
rect 688 161 697 195
rect 697 161 731 195
rect 731 161 740 195
rect 688 144 740 161
<< metal2 >>
rect 0 1149 884 1155
rect 0 1148 382 1149
rect 0 1096 140 1148
rect 192 1096 382 1148
rect 0 1084 382 1096
rect 0 1032 140 1084
rect 192 1032 382 1084
rect 0 1020 382 1032
rect 0 968 140 1020
rect 192 968 382 1020
rect 0 956 382 968
rect 0 904 140 956
rect 192 905 382 956
rect 498 1097 688 1149
rect 740 1097 884 1149
rect 498 1085 884 1097
rect 498 1033 688 1085
rect 740 1033 884 1085
rect 498 1021 884 1033
rect 498 969 688 1021
rect 740 969 884 1021
rect 498 957 884 969
rect 498 905 688 957
rect 740 905 884 957
rect 192 904 884 905
rect 0 898 884 904
rect 0 864 884 870
rect 0 428 228 864
rect 344 428 536 864
rect 652 428 884 864
rect 0 422 884 428
rect 0 388 884 394
rect 0 336 140 388
rect 192 336 688 388
rect 740 336 884 388
rect 0 324 884 336
rect 0 272 140 324
rect 192 272 688 324
rect 740 272 884 324
rect 0 260 884 272
rect 0 208 140 260
rect 192 208 688 260
rect 740 208 884 260
rect 0 196 884 208
rect 0 144 140 196
rect 192 144 688 196
rect 740 144 884 196
rect 0 138 884 144
<< labels >>
flabel comment s 278 681 278 681 0 FreeSans 300 0 0 0 D
flabel comment s 737 681 737 681 0 FreeSans 300 0 0 0 S
flabel comment s 432 681 432 681 0 FreeSans 300 0 0 0 S
flabel comment s 158 681 158 681 0 FreeSans 300 180 0 0 S
flabel comment s 586 681 586 681 0 FreeSans 300 0 0 0 D
flabel metal1 s 414 50 500 75 0 FreeSans 200 180 0 0 GATE
port 2 nsew
flabel metal2 s 233 599 309 624 0 FreeSans 200 0 0 0 DRAIN
port 3 nsew
flabel metal2 s 0 1055 76 1080 0 FreeSans 200 0 0 0 SOURCE
port 4 nsew
flabel mvpdiff s 52 722 52 722 0 FreeSans 700 270 0 0 Bulk
<< properties >>
string GDS_END 10042372
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10013450
<< end >>
