magic
tech sky130A
magscale 1 2
timestamp 1746986264
<< obsli1 >>
rect -1140 7100 1290 7182
rect -1140 -1100 -1058 7100
rect -962 9 -896 5991
rect 8 43 142 5957
rect 1046 9 1112 5991
rect -296 -857 460 -643
rect 1208 -1100 1290 7100
rect -1140 -1182 1290 -1100
<< obsm1 >>
rect -1140 7100 1290 7182
rect -1140 -1100 -1058 7100
rect -958 19 -900 5981
rect 10 55 140 5945
rect 1050 19 1108 5981
rect -296 -857 460 -643
rect 1208 -1100 1290 7100
rect -1140 -1182 1290 -1100
<< obsm2 >>
rect 11 57 139 5945
rect -296 -857 460 -643
<< properties >>
string FIXED_BBOX 0 0 2430 8364
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7579874
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 7459866
<< end >>
