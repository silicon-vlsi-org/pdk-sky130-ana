* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* ./models_diodes.spice created from ./models.spice
*
**********************************
******************************************************************
******************************************************************
*  *****************************************************
*  04/05/2021 Usman Suriono
*      Why     : New infrastructure of diode models
*      What    : Converted from sky130_fd_pr__model__parasitic__diode_ps2dn_n20zvtvh1defet model
*                Added estimated breakdown Corners
*
*  *****************************************************
*
*  Deep Nwell Extended Drain to Substrate Model
*  Based on the layout 20V Nmos Zero VT device
*  -----------------------------------------------------

.subckt  sky130_fd_pr__model__parasitic__diode_ps2dn__extended_drain a c mult=1
+ area=1 perim=1
+ 
.param  sky130_fd_pr__nfet_20v0_zvt_cjdnwpsubjunction_mult = 7.0510e-01
+ sky130_fd_pr__nfet_20v0_zvt_mjdnwpsubjunction_mult = 1.6541
+ sky130_fd_pr__nfet_20v0_zvt_pbdnwpsubjunction_mult = 1.4206
+ sky130_fd_pr__nfet_20v0_zvt_vb = {30.0/(1+0.2*(sw_func_dnw_sub_cj-1))}


Dsky130_fd_pr__model__parasitic__diode_ps2dn__extended_drain a c sky130_fd_pr__model__parasitic__diode_ps2dn_diode area = {area} pj = {perim}


.model sky130_fd_pr__model__parasitic__diode_ps2dn_diode d 
+ level = 3
*
*PARAMETERS TO MAKE MODEL INTO CADFLOW
*
+ tlevc = 1
+ area = 1e12
*
*JUNCTION CAPACITANCE PARAMETERS
*
+ cj = {1.176E-04*1e-12*sw_func_dnw_sub_cj}
+ mj = {0.56056*sky130_fd_pr__nfet_20v0_zvt_mjdnwpsubjunction_mult}
+ pb = {0.21294*sky130_fd_pr__nfet_20v0_zvt_pbdnwpsubjunction_mult}
+ cjsw = {8.1380e-010*sky130_fd_pr__nfet_20v0_zvt_cjdnwpsubjunction_mult*1e-6*sw_func_dnw_sub_cj}
+ mjsw = {0.18742*sky130_fd_pr__nfet_20v0_zvt_mjdnwpsubjunction_mult}
+ php = {0.21294*sky130_fd_pr__nfet_20v0_zvt_pbdnwpsubjunction_mult}
+ cta = 0.0031223
+ ctp = 0.0014703
+ tpb = 0.0016859
+ tphp = 0.0016859
*
*DIODE IV PARAMETERS
*
+ js = 6.1049e-017
+ jsw = 8.1115e-016
+ n = 0.9891
+ rs = {900*1e-12}
+ ik = {2.08e-009/1e-12}
+ ikr = 0
******set to 40V so design can evaluate circuits using up to 36V
+ bv = {sky130_fd_pr__nfet_20v0_zvt_vb}
+ ibv = 0.00106
+ trs = 0
+ eg = 1.17
+ xti = 1.0
+ tref = 30
*
*DEFAULT PARAMETERS
*
+ tcv = 0
+ gap1 = 0.000473
+ gap2 = 1110
+ ttt1 = 0
+ ttt2 = 0
+ tm1 = 0
+ tm2 = 0
+ lm = 0
+ lp = 0
+ wm = 0
+ wp = 0
+ xm = 0
+ xoi = 10000
+ xom = 10000
+ xp = 0
+ xw = 0

.ends sky130_fd_pr__model__parasitic__diode_ps2dn__extended_drain
******************************************************************
******************************************************************
*  *****************************************************
*  02/16/2021 Usman Suriono
*      Why     : New infrastructure of diode models
*      What    : Converted from dnwdiode_psub model
*                Added estimated breakdown Corners.
*
*  *****************************************************
*
*  Deep Nwell to Substrate Model
*  -----------------------------------------------------


.subckt  sky130_fd_pr__model__parasitic__diode_ps2dn a c mult=1
+ area=1 perim=1

Dsky130_fd_pr__model__parasitic__diode_ps2dn a c sky130_fd_pr__model__parasitic__diode_ps2dn_diode area = {area} pj = {perim}


.model sky130_fd_pr__model__parasitic__diode_ps2dn_diode d 

+ level = 3
*
*PARAMETERS TO MAKE MODEL INTO CADFLOW
*
+ tlevc = 1
+ area = 1e12
*
*JUNCTION CAPACITANCE PARAMETERS
*
+ cj = {sw_dnw_sub_cj*1e-12}
+ mj = 0.49
+ pb = 0.5348
+ cjsw = {8.1664e-010*1e-6*sw_func_dnw_sub_cj}
+ mjsw = 0.20024
+ php = 0.5348
+ cta = 0.0016157
+ ctp = 0.0008
+ tpb = 0.0025003
+ tphp = 0.001675
*
*DIODE IV PARAMETERS
*
+ js = 6.1049e-017
+ jsw = 8.1115e-016
+ n = 1.0791
+ rs = {900*1e-12}
+ ik = {2.08e-009/1e-12}
+ ikr = {0/1e-12}
+ bv = {16.95/(1+0.2*(sw_func_dnw_sub_cj-1))}
+ ibv = 0.00106
+ trs = 0
+ eg = 1.17
+ xti = 1.0
+ tref = 30
*
*DEFAULT PARAMETERS
*
+ tcv = 0
+ gap1 = 0.000473
+ gap2 = 1110
+ ttt1 = 0
+ ttt2 = 0
+ tm1 = 0
+ tm2 = 0
+ lm = 0
+ lp = 0
+ wm = 0
+ wp = 0
+ xm = 0
+ xoi = 10000
+ xom = 10000
+ xp = 0
+ xw = 0

.ends sky130_fd_pr__model__parasitic__diode_ps2dn
******************************************************************
******************************************************************
*  *****************************************************
*  04/05/2021 Usman Suriono
*      Why     : New model structure
*      What    : Converted from dnwdiode_pw_defet models
*                Added estimated Corner breakdown
*
*  *****************************************************
*
*  Isolated Pwell to Nwell Diode for Extended Drain Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__model__parasitic__diode_pw2dn_defet a c mult=1
+ area=1 perim=1

Dsky130_fd_pr__model__parasitic__diode_pw2dn_defet a c diodeint area = {area} pj = {perim}


.model diodeint d 
+ level = 3
*
*PARAMETERS TO MAKE MODEL INTO CADFLOW
*
+ tlevc = 1
+ area = 1e12
*
*JUNCTION CAPACITANCE PARAMETERS
*
+ cj = {sw_pw_dnw_cj*1e-12*7.5058e-01}
+ mj = {0.63982*8.3390e-01}
+ pb = {0.58758*1.0204e+00}
+ cjsw = {3.743e-010*1e-6*sw_func_pw_dnw_cj*7.5058e-01}
+ mjsw = {0.80357*8.3390e-01}
+ php = {0.2500*1.0204e+00}
+ cta = 0.0016157
+ ctp = 0.0008
+ tpb = 0.0010003
+ tphp = 0.000675
*
*DIODE IV PARAMETERS
*
+ minr = 1e-3
+ js = 1.4693e-017
+ jsw = 7.41e-018
+ n = 1.0791
+ rs = {900*1e-12}
+ ik = {2.08e-009/1e-12}
+ ikr = {0/1e-12}
******set to 40V so design can evaluate circuits using up to 36V
+ bv = {26/(1+0.3*(sw_func_pw_dnw_cj-1))}
+ ibv = 0.00106
+ trs = 0
+ xti = 3.0
+ eg = 1.50
+ tref = 30
*
*DEFAULT PARAMETERS
*
+ tcv = 0
+ gap1 = 0.000473
+ gap2 = 1110
+ ttt1 = 0
+ ttt2 = 0
+ tm1 = 0
+ tm2 = 0
+ lm = 0
+ lp = 0
+ wm = 0
+ wp = 0
+ xm = 0
+ xoi = 10000
+ xom = 10000
+ xp = 0
+ xw = 0

.ends sky130_fd_pr__model__parasitic__diode_pw2dn_defet
******************************************************************
******************************************************************
*  *****************************************************
*  02/19/2021 Usman Suriono
*      Why     : New model structure
*      What    : Converted from dnwdiode_pw model
*                Add estimated BV Corners
*
*  *****************************************************
*
*  Isolated Pwell to Nwell Diode Model
*  -----------------------------------------------------


.subckt  sky130_fd_pr__model__parasitic__diode_pw2dn a c mult=1
+ area=1 perim=1

Dsky130_fd_pr__model__parasitic__diode_pw2dn a c diodeint area = {area} pj = {perim}


.model diodeint d 
+ level = 3
*
*PARAMETERS TO MAKE MODEL INTO CADFLOW
*
+ tlevc = 1
+ area = 1e12
*
*JUNCTION CAPACITANCE PARAMETERS
*
+ cj = {sw_pw_dnw_cj*1e-12}
+ mj = 0.33982
+ pb = 0.58758
+ cjsw = {3.743e-010*1e-6*sw_func_pw_dnw_cj}
+ mjsw = 0.23357
+ php = 0.5348
+ cta = 0.0016157
+ ctp = 0.0008
+ tpb = 0.0025003
+ tphp = 0.001675
*
*DIODE IV PARAMETERS
*
+ js = 1.4693e-017
+ jsw = 7.41e-018
+ n = 1.0791
+ rs = {900*1e-12}
+ ik = {2.08e-009/1e-12}
+ ikr = {0/1e-12}
+ bv = {16.38/(1+0.3*(sw_func_pw_dnw_cj-1))}
+ ibv = 0.00106
+ trs = 0
+ eg = 1.17
+ xti = 3.0
+ tref = 30
*
*DEFAULT PARAMETERS
*
+ tcv = 0
+ gap1 = 0.000473
+ gap2 = 1110
+ ttt1 = 0
+ ttt2 = 0
+ tm1 = 0
+ tm2 = 0
+ lm = 0
+ lp = 0
+ wm = 0
+ wp = 0
+ xm = 0
+ xoi = 10000
+ xom = 10000
+ xp = 0
+ xw = 0

.ends sky130_fd_pr__model__parasitic__diode_pw2dn
******************************************************************
******************************************************************
*  *****************************************************
*  12/16/2020 Usman Suriono
*      Why     : New infrastructure of diode models
*      What    : Converted from ndiode_defet model
*                This model is identical to sky130_fd_pr__diode_pw2nd_05v5 except for higher "pb" parameter
*
*  *****************************************************
*
*  Junction diode of S/B of Nmos 20V VHV DE for Extend Drain Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__diode_pw2nd_05v5_defet a c mult=1
+ area=1 perim=1

Dsky130_fd_pr__diode_pw2nd_05v5_defet a c diodeint area = {area} pj = {perim}


.model diodeint d minr = 0.001
+ level = 3
*
*PARAMETERS TO MAKE MODEL INTO CADFLOW
*
+ tlevc = 1
+ area = 1e12
*
*JUNCTION CAPACITANCE PARAMETERS
*
+ cj = {sw_nsd_pw_cj*1e-12}
+ mj = 0.44
+ pb = {0.729*2.7281}
+ cjsw = {3.6001e-011*1e-6*sw_func_nsd_pw_cj}
+ mjsw = 0.0009
+ php = 0.2
+ cta = 0.000792
+ ctp = 1e-005
+ tpb = 0.0012287
+ tphp = 0
*
*DIODE IV PARAMETERS
*
+ js = 2.75e-015
+ jsw = 6e-016
+ n = 1.2928
+ rs = {981*1e-12}
+ ik = {1.3e-009/1e-12}
+ ikr = {0/1e-12}
+ bv = {11.7/sw_func_nsd_pw_cj}
+ ibv = 0.00106
+ trs = 0
+ eg = 1.05
+ xti = 2
+ tref = 30
*
*DEFAULT PARAMETERS
*
+ tcv = 0
+ gap1 = 0.000473
+ gap2 = 1110
+ ttt1 = 0
+ ttt2 = 0
+ tm1 = 0
+ tm2 = 0
+ lm = 0
+ lp = 0
+ wm = 0
+ wp = 0
+ xm = 0
+ xoi = 10000
+ xom = 10000
+ xp = 0
+ xw = 0

.ends sky130_fd_pr__diode_pw2nd_05v5_defet
******************************************************************
******************************************************************
*  *****************************************************
*  03/06/2021 Usman Suriono
*      Why     : New model structure
*      What    : Converted from xesd_ndiode_h_100 model
*                Added estimated Corners for breakdown
*
*  *****************************************************
*
*  ESD NPlus to Pwell Diode Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__diode_pw2nd_05v5_esd c0 c1 mult=1
+ area=1 perim=1
xd1 a1 c1 sky130_fd_pr__diode_pw2nd_05v5 area = {area*1.54} perim = {perim} rs_int = {0*1e-12}
Rsky130_fd_pr__diode_pw2nd_05v5_esd c0 a1 r = 1.1101


.ends sky130_fd_pr__diode_pw2nd_05v5_esd

******************************************************************
******************************************************************
*  *****************************************************
*  03/06/2021 Usman Suriono
*      Why     : New model structure
*      What    : Converted from xesd_ndiode_h_100 model
*                Added estimated Corners for breakdown
*
*  *****************************************************
*
*  ESD NPlus to Pwell Diode Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__diode_pw2nd_05v5_esd_v5 c0 c1 mult=1
+ area=1 perim=1
xd1 a1 c1 sky130_fd_pr__diode_pw2nd_11v0 area = {area*1.54} perim = {perim} rs_int = {0*1e-12}
Rsky130_fd_pr__diode_pw2nd_05v5_esd_v5 c0 a1 r = 1.1101


.ends sky130_fd_pr__diode_pw2nd_05v5_esd_v5

******************************************************************
******************************************************************
*  *****************************************************
*  11/10/2020 Usman Suriono
*      Why     : New model structure
*      What    : Converted from ndiode_lvt model
*                Added estimated Corner for breakdwon
*
*  *****************************************************
*
*  NPlus to Pwell Low VT Diode Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__diode_pw2nd_05v5_lvt a c mult=1
+ area=1 perim=1

Dsky130_fd_pr__diode_pw2nd_05v5_lvt a c diodeint area = {area} pj = {perim}


.model diodeint d 
+ level = 3
*
*PARAMETERS TO MAKE MODEL INTO CADFLOW
*
+ tlevc = 1
+ area = 1e12
*
*JUNCTION CAPACITANCE PARAMETERS
*
+ cj = {1.210E-03*1e-12*sw_func_nsd_pw_cj}
+ mj = 0.42197
+ pb = 0.7477
+ cjsw = {3.6224e-011*1e-6*sw_func_nsd_pw_cj}
+ mjsw = 0.001
+ php = 0.1
+ cta = 0.000792
+ ctp = 1e-005
+ tpb = 0.0012287
+ tphp = 0
*
*DIODE IV PARAMETERS
*
+ js = 2.75e-015
+ jsw = 6e-016
+ n = 1.2928
+ rs = {981*1e-12}
+ ik = {1.3e-009/1e-12}
+ ikr = {0/1e-12}
+ bv = {11.9/sw_func_nsd_pw_cj}
+ ibv = 0.00106
+ trs = 0
+ eg = 1.05
+ xti = 2
+ tref = 30
*
*DEFAULT PARAMETERS
*
+ tcv = 0
+ gap1 = 0.000473
+ gap2 = 1110
+ ttt1 = 0
+ ttt2 = 0
+ tm1 = 0
+ tm2 = 0
+ lm = 0
+ lp = 0
+ wm = 0
+ wp = 0
+ xm = 0
+ xoi = 10000
+ xom = 10000
+ xp = 0
+ xw = 0

.ends sky130_fd_pr__diode_pw2nd_05v5_lvt
******************************************************************
******************************************************************
*  *****************************************************
*  11/10/2020 Usman Suriono
*      Why     : New model structure
*      What    : Converted from ndiode_native model
*
*  *****************************************************
*
*  NPlus to Pwell Native VT Diode Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__diode_pw2nd_05v5_nvt a c mult=1
+ area=1 perim=1

Dsky130_fd_pr__diode_pw2nd_05v5_nvt a c diodeint area = {area} pj = {perim}


.model diodeint d 
+ level = 3
*
*PARAMETERS TO MAKE MODEL INTO CADFLOW
*
+ tlevc = 1
+ area = 1e12
*
*JUNCTION CAPACITANCE PARAMETERS
*
+ cj = {8.310E-04*1e-12*sw_func_nsd_pw_cj}
+ mj = 0.28329
+ pb = 0.66345
+ cjsw = {8.5152e-011*1e-6*sw_func_nsd_pw_cj}
+ mjsw = 0.057926
+ php = 1
+ cta = 0.00083
+ ctp = 0
+ tpb = 0.0019685
+ tphp = 0.001
*
*DIODE IV PARAMETERS
*
+ js = 4.2966e-016
+ jsw = 8.04e-016
+ n = 1.5764
+ rs = {600*1e-12}
+ ik = {4.76e-008/1e-12}
+ ikr = {0/1e-12}
+ bv = {12.69/sw_func_nsd_pw_cj}
+ ibv = 0.00106
+ trs = 0
+ eg = 1.05
+ xti = 0
+ tref = 30
*
*DEFAULT PARAMETERS
*
+ tcv = 0
+ gap1 = 0.000473
+ gap2 = 1110
+ ttt1 = 0
+ ttt2 = 0
+ tm1 = 0
+ tm2 = 0
+ lm = 0
+ lp = 0
+ wm = 0
+ wp = 0
+ xm = 0
+ xoi = 10000
+ xom = 10000
+ xp = 0
+ xw = 0

.ends sky130_fd_pr__diode_pw2nd_05v5_nvt
******************************************************************
******************************************************************
*  *****************************************************
*  11/10/2020 Usman Suriono
*      Why     : New model structure
*      What    : Converted from ndiode model
*                Added estimated Corners for breakdown
*
*  *****************************************************
*
*  NPlus to Pwell normal sky130_fd_pr__nfet_01v8 VT Diode Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__diode_pw2nd_05v5 a c mult=1
+ area=1 perim=1 
.param  rs_int = {981*1e-12}

Dsky130_fd_pr__diode_pw2nd_05v5 a c ndiode area = {area} pj = {perim}


.model ndiode d 
+ level = 3
*
*PARAMETERS TO MAKE MODEL INTO CADFLOW
*
+ tlevc = 1
+ area = 1e12
*
*JUNCTION CAPACITANCE PARAMETERS
*
+ cj = {sw_nsd_pw_cj*1e-12}
+ mj = 0.44
+ pb = 0.729
+ cjsw = {3.6001e-011*1e-6*sw_func_nsd_pw_cj}
+ mjsw = 0.0009
+ php = 0.2
+ cta = 0.000792
+ ctp = 1e-005
+ tpb = 0.0012287
+ tphp = 0
*
*DIODE IV PARAMETERS
*
+ js = 2.75e-015
+ jsw = 6e-016
+ n = 1.2928
+ rs = {rs_int}
+ ik = {1.3e-009/1e-12}
+ ikr = 0
+ bv = {11.7/sw_func_nsd_pw_cj}
+ ibv = 0.00106
+ trs = 0
+ eg = 1.05
+ xti = 2
+ tref = 30
*
*DEFAULT PARAMETERS
*
+ tcv = 0
+ gap1 = 0.000473
+ gap2 = 1110
+ ttt1 = 0
+ ttt2 = 0
+ tm1 = 0
+ tm2 = 0
+ lm = 0
+ lp = 0
+ wm = 0
+ wp = 0
+ xm = 0
+ xoi = 10000
+ xom = 10000
+ xp = 0
+ xw = 0

.ends sky130_fd_pr__diode_pw2nd_05v5
******************************************************************
******************************************************************
*  *****************************************************
*  11/10/2020 Usman Suriono
*      Why     : New model structure
*      What    : Converted from ndiode_h models
*                Added estimated Corner for breakdown
*
*  *****************************************************
*
*  NPlus to Pwell 5V Diode Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__diode_pw2nd_11v0 a c mult=1
+ area=1 perim=1 
.param  rs_int = {981*1e-12}

Dsky130_fd_pr__diode_pw2nd_11v0 a c ndiode_h area = {area} pj = {perim}


.model ndiode_h d 
+ level = 3
*
*PARAMETERS TO MAKE MODEL INTO CADFLOW
*
+ tlevc = 1
+ area = 1e12
*
*JUNCTION CAPACITANCE PARAMETERS
*
+ cj = {0.0008512*1e-12*sw_func_nsd_pw_cj}
+ mj = 0.295
+ pb = 0.72468
+ cjsw = {8.5204e-011*1e-6*sw_func_nsd_pw_cj}
+ mjsw = 0.037586
+ php = 0.29067
+ cta = 0.00067434
+ ctp = 0.0002493
+ tpb = 0.001344
+ tphp = 0.00099005
*
*DIODE IV PARAMETERS
*
+ js = 3.75e-016
+ jsw = 5.84e-017
+ n = 1.0773
+ rs = {rs_int}
+ ik = {1.3e-009/1e-12}
+ ikr = {0/1e-12}
+ bv = {12.636/sw_func_nsd_pw_cj}
+ ibv = 0.00106
+ trs = 0
+ eg = 0.92
+ xti = 0.76
+ tref = 30
*
*DEFAULT PARAMETERS
*
+ tcv = 0
+ gap1 = 0.000473
+ gap2 = 1110
+ ttt1 = 0
+ ttt2 = 0
+ tm1 = 0
+ tm2 = 0
+ lm = 0
+ lp = 0
+ wm = 0
+ wp = 0
+ xm = 0
+ xoi = 10000
+ xom = 10000
+ xp = 0
+ xw = 0

.ends sky130_fd_pr__diode_pw2nd_11v0
******************************************************************
******************************************************************
*  *****************************************************
*  02/13/2021 Usman Suriono
*      Why     : New model structure
*      What    : Converted from nwdiode model
*                Add estimated BV Corners
*
*  *****************************************************
*
*  Nwell to isolated Pwell Diode Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__model__parasitic__diode_pd2nw a c mult=1
+ area=1 perim=1

Dsky130_fd_pr__model__parasitic__diode_pd2nw a c diodeint area = {area} pj = {perim}


.model diodeint d 
+ level = 3
*
*PARAMETERS TO MAKE MODEL INTO CADFLOW
*
+ tlevc = 1
+ area = 1e12
*
*JUNCTION CAPACITANCE PARAMETERS
*
+ cj = {sw_nw_pw_cj*1e-12}
+ mj = 0.4509
+ pb = 0.5348
+ cjsw = {5.822e-010*1e-6*sw_func_nw_pw_cj}
+ mjsw = 0.2433
+ php = 0.5348
+ cta = 0.00165
+ ctp = 0.0008
+ tpb = 0.0022563
+ tphp = 0.00165
*
*DIODE IV PARAMETERS
*
+ js = 4.21e-018
+ jsw = 4.94e-018
+ n = 1.0791
+ rs = {900*1e-12}
+ ik = {2.08e-009/1e-12}
+ ikr = {0/1e-12}
+ bv = {16.848/sw_func_nw_pw_cj}
+ ibv = 0.00106
+ trs = 0
+ eg = 1.17
+ xti = 5.2
+ tref = 30
*
*DEFAULT PARAMETERS
*
+ tcv = 0
+ gap1 = 0.000473
+ gap2 = 1110
+ ttt1 = 0
+ ttt2 = 0
+ tm1 = 0
+ tm2 = 0
+ lm = 0
+ lp = 0
+ wm = 0
+ wp = 0
+ xm = 0
+ xoi = 10000
+ xom = 10000
+ xp = 0
+ xw = 0

.ends sky130_fd_pr__model__parasitic__diode_pd2nw
******************************************************************
******************************************************************
*  *****************************************************
*  02/17/2021 Usman Suriono
*      Why     : New model structure
*      What    : Converted from dnwdiode_psub model
*                Added estimated Corner for breakdwon
*                The junction cap follows lower doping, correlated to PSD-NW
*
*  *****************************************************
*
*  Photo Diode Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__photodiode a c mult=1
+ area=1 perim=1

Dsky130_fd_pr__photodiode a c diodeint area = {area} pj = {perim}


.model diodeint d 
+ level = 3
*
*PARAMETERS TO MAKE MODEL INTO CADFLOW
*
+ tlevc = 1
+ area = 1e12
*
*JUNCTION CAPACITANCE PARAMETERS
*
+ cj = {7.8544e-005*1e-12*sw_func_psd_nw_cj}
+ mj = 0.49
+ pb = 0.5348
+ cjsw = {8.1664e-010*1e-6*sw_func_psd_nw_cj}
+ mjsw = 0.20024
+ php = 0.5348
+ cta = 0.0016157
+ ctp = 0.0008
+ tpb = 0.0025003
+ tphp = 0.001675
*
*DIODE IV PARAMETERS
*
+ js = 6.1049e-017
+ jsw = 8.1115e-016
+ n = 1.0791
+ rs = {900*1e-12}
+ ik = {2.08e-009/1e-12}
+ ikr = {0/1e-12}
+ bv = {16.95/sw_func_psd_nw_cj}
+ ibv = 0.00106
+ trs = 0
+ eg = 1.17
+ xti = 1.0
+ tref = 30
*
*DEFAULT PARAMETERS
*
+ tcv = 0
+ gap1 = 0.000473
+ gap2 = 1110
+ ttt1 = 0
+ ttt2 = 0
+ tm1 = 0
+ tm2 = 0
+ lm = 0
+ lp = 0
+ wm = 0
+ wp = 0
+ xm = 0
+ xoi = 10000
+ xom = 10000
+ xp = 0
+ xw = 0

.ends sky130_fd_pr__photodiode
******************************************************************
******************************************************************
*  *****************************************************
*  03/06/2021 Usman Suriono
*      Why     : New model structure
*      What    : Converted from xesd_ndiode_h_100 model
*                Added estimated Corners for breakdown
*
*  *****************************************************
*
*  ESD NPlus to Pwell Diode Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__diode_pd2nw_05v5_esd c0 c1 mult=1
+ area=1 perim=1
xd1 a1 c1 sky130_fd_pr__diode_pd2nw_05v5 area = {area*1.54} perim = {perim} rs_int = {0*1e-12}
Rsky130_fd_pr__diode_pd2nw_05v5_esd c0 a1 r = 1.1101


.ends sky130_fd_pr__diode_pd2nw_05v5_esd

******************************************************************
******************************************************************
*  *****************************************************
*  03/06/2021 Usman Suriono
*      Why     : New model structure
*      What    : Converted from xesd_ndiode_h_100 model
*                Added estimated Corners for breakdown
*
*  *****************************************************
*
*  ESD NPlus to Pwell Diode Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__diode_pd2nw_05v5_esd_v5 c0 c1 mult=1
+ area=1 perim=1
xd1 a1 c1 sky130_fd_pr__diode_pd2nw_11v0 area = {area*1.54} perim = {perim} rs_int = {0*1e-12}
Rsky130_fd_pr__diode_pd2nw_05v5_esd_v5 c0 a1 r = 1.1101


.ends sky130_fd_pr__diode_pd2nw_05v5_esd_v5

******************************************************************
******************************************************************
*  *****************************************************
*  02/13/2021 Usman Suriono
*      Why     : New model structure
*      What    : Converted from pdiode_hvt model
*                Add estimated BV Corners
*
*  *****************************************************
*
*  PPlus to Nwell Pmos High VT Diode Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__diode_pd2nw_05v5_hvt a c mult=1
+ area=1 perim=1


Dsky130_fd_pr__diode_pd2nw_05v5_hvt a c diodeint area = {area} pj = {perim}



.model diodeint d 
+ level = 3
*
*PARAMETERS TO MAKE MODEL INTO CADFLOW
*
+ tlevc = 1
+ area = 1e12
*
*JUNCTION CAPACITANCE PARAMETERS
*
+ cj = {7.433E-04*1e-12*sw_func_psd_nw_cj}
+ mj = 0.34629
+ pb = 0.6587
+ cjsw = {9.2435e-011*1e-6*sw_func_psd_nw_cj}
+ mjsw = 0.26859
+ php = 0.7418
+ cta = 0.0012407
+ ctp = 0
+ tpb = 0.0019551
+ tphp = 0.00014242
*
*DIODE IV PARAMETERS
*
+ js = 2.17e-017
+ jsw = 8.2e-016
+ n = 1.2556
+ rs = {600*1e-12}
+ ik = {4.76e-008/1e-12}
+ ikr = {0/1e-12}
+ bv = {12.8/sw_func_psd_nw_cj}
+ ibv = 0.00106
+ trs = 0
+ eg = 1.05
+ xti = 2.0
+ tref = 30
*
*DEFAULT PARAMETERS
*
+ tcv = 0
+ gap1 = 0.000473
+ gap2 = 1110
+ ttt1 = 0
+ ttt2 = 0
+ tm1 = 0
+ tm2 = 0
+ lm = 0
+ lp = 0
+ wm = 0
+ wp = 0
+ xm = 0
+ xoi = 10000
+ xom = 10000
+ xp = 0
+ xw = 0

.ends sky130_fd_pr__diode_pd2nw_05v5_hvt
******************************************************************
******************************************************************
*  *****************************************************
*  12/03/2020 Usman Suriono
*      Why     : New model structure
*      What    : Converted from pdiode_lvt model
*                Add estimated BV Corners
*
*  *****************************************************
*
*  PPlus to Nwell Pmos Low VT Diode Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__diode_pd2nw_05v5_lvt a c mult=1
+ area=1 perim=1


Dsky130_fd_pr__diode_pd2nw_05v5_lvt a c  diodeint area = {area} pj = {perim}


.model diodeint d 
+ level = 3
*
*PARAMETERS TO MAKE MODEL INTO CADFLOW
*
+ tlevc = 1
+ area = 1e12
*
*JUNCTION CAPACITANCE PARAMETERS
*
+ cj = {7.682E-04*1e-12*sw_func_psd_nw_cj}
+ mj = 0.3362
+ pb = 0.6587
+ cjsw = {9.152e-011*1e-6*sw_func_psd_nw_cj}
+ mjsw = 0.2659
+ php = 0.7418
+ cta = 0.0012407
+ ctp = 0.00037357
+ tpb = 0.001671
+ tphp = 0.001246
*
*DIODE IV PARAMETERS
*
+ js = 2.1483e-017
+ jsw = 1.447e-16
+ n = 1.3632
+ rs = {600*1e-12}
+ ik = {4.76e-008/1e-12}
+ ikr = {0/1e-12}
+ bv = {12.69/sw_func_psd_nw_cj}
+ ibv = 0.00106
+ trs = 0
+ eg = 1.05
+ xti = 5.2
+ tref = 30
*
*DEFAULT PARAMETERS
*
+ tcv = 0
+ gap1 = 0.000473
+ gap2 = 1110
+ ttt1 = 0
+ ttt2 = 0
+ tm1 = 0
+ tm2 = 0
+ lm = 0
+ lp = 0
+ wm = 0
+ wp = 0
+ xm = 0
+ xoi = 10000
+ xom = 10000
+ xp = 0
+ xw = 0

.ends sky130_fd_pr__diode_pd2nw_05v5_lvt
******************************************************************
******************************************************************
*  *****************************************************
*  12/03/2020 Usman Suriono
*      Why     : New model structure
*      What    : Converted from pdiode model
*                Add estimated BV Corners
*
*  *****************************************************
*
*  PPlus to Nwell normal Pmos VT Diode Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__diode_pd2nw_05v5 a c mult=1
+ area=1 perim=1 
.param  rs_int = {600*1e-12}

Dsky130_fd_pr__diode_pd2nw_05v5 a c pdiode area = {area} pj = {perim}



.model pdiode d 
+ level = 3
*
*PARAMETERS TO MAKE MODEL INTO CADFLOW
*
+ tlevc = 1
+ area = 1e12
*
*JUNCTION CAPACITANCE PARAMETERS
*
+ cj = {sw_psd_nw_cj*1e-12}
+ mj = 0.34629
+ pb = 0.6587
+ cjsw = {9.88e-011*1e-6*sw_func_psd_nw_cj}
+ mjsw = 0.29781
+ php = 0.7418
+ cta = 0.0012407
+ ctp = 0.00037357
+ tpb = 0.0020386
+ tphp = 0.001246
*
*DIODE IV PARAMETERS
*
+ js = 2.1483e-017
+ jsw = 8.04e-016
+ n = 1.3632
+ rs = {rs_int}
+ ik = {4.76e-008/1e-12}
+ ikr = 0
+ bv = {12.69/sw_func_psd_nw_cj}
+ ibv = 0.00106
+ trs = 0
+ eg = 1.05
+ xti = 5.2
+ tref = 30
*
*DEFAULT PARAMETERS
*
+ tcv = 0
+ gap1 = 0.000473
+ gap2 = 1110
+ ttt1 = 0
+ ttt2 = 0
+ tm1 = 0
+ tm2 = 0
+ lm = 0
+ lp = 0
+ wm = 0
+ wp = 0
+ xm = 0
+ xoi = 10000
+ xom = 10000
+ xp = 0
+ xw = 0

.ends sky130_fd_pr__diode_pd2nw_05v5
******************************************************************
******************************************************************
*  *****************************************************
*  02/13/2021 Usman Suriono
*      Why     : New model structure
*      What    : Converted from pdiode_h model
*                Add estimated BV Corners
*
*  *****************************************************
*
*  PPlus to Nwell 5V Diode Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__diode_pd2nw_11v0 a c mult=1
+ area=1 perim=1 
.param  rs_int = {600*1e-12}

Dsky130_fd_pr__diode_pd2nw_11v0 a c pdiode_h area = {area} pj = {perim}


.model pdiode_h d 
+ level = 3
*
*PARAMETERS TO MAKE MODEL INTO CADFLOW
*
+ tlevc = 1
+ area = 1e12
*
*JUNCTION CAPACITANCE PARAMETERS
*
+ cj = {0.00077547*1e-12*sw_func_psd_nw_cj}
+ mj = 0.33956
+ pb = 0.6587
+ cjsw = {9.8717e-011*1e-6*sw_func_psd_nw_cj}
+ mjsw = 0.24676
+ php = 1
+ cta = 0.00096
+ ctp = 3e-005
+ tpb = 0.001671
+ tphp = 0
*
*DIODE IV PARAMETERS
*
+ js = 2.1483e-017
+ jsw = 4.02e-018
+ n = 1.3632
+ rs = {rs_int}
+ ik = {4.76e-008/1e-12}
+ ikr = 0
+ bv = {12.69/sw_func_psd_nw_cj}
+ ibv = 0.00106
+ trs = 0
+ eg = 1.05
+ xti = 10
+ tref = 30
*
*DEFAULT PARAMETERS
*
+ tcv = 0
+ gap1 = 0.000473
+ gap2 = 1110
+ ttt1 = 0
+ ttt2 = 0
+ tm1 = 0
+ tm2 = 0
+ lm = 0
+ lp = 0
+ wm = 0
+ wp = 0
+ xm = 0
+ xoi = 10000
+ xom = 10000
+ xp = 0
+ xw = 0

.ends sky130_fd_pr__diode_pd2nw_11v0
