magic
tech sky130A
magscale 1 2
timestamp 1746986264
<< locali >>
rect 167 1160 179 1194
rect 213 1160 251 1194
rect 285 1160 323 1194
rect 357 1160 369 1194
rect 48 1020 82 1058
rect 48 948 82 986
rect 48 876 82 914
rect 48 804 82 842
rect 48 732 82 770
rect 48 660 82 698
rect 48 588 82 626
rect 48 516 82 554
rect 48 444 82 482
rect 48 372 82 410
rect 48 300 82 338
rect 48 228 82 266
rect 48 122 82 194
rect 454 1020 488 1058
rect 454 948 488 986
rect 454 876 488 914
rect 454 804 488 842
rect 454 732 488 770
rect 454 660 488 698
rect 454 588 488 626
rect 454 516 488 554
rect 454 444 488 482
rect 454 372 488 410
rect 454 300 488 338
rect 454 228 488 266
rect 454 122 488 194
rect 167 20 179 54
rect 213 20 251 54
rect 285 20 323 54
rect 357 20 369 54
<< viali >>
rect 179 1160 213 1194
rect 251 1160 285 1194
rect 323 1160 357 1194
rect 48 1058 82 1092
rect 48 986 82 1020
rect 48 914 82 948
rect 48 842 82 876
rect 48 770 82 804
rect 48 698 82 732
rect 48 626 82 660
rect 48 554 82 588
rect 48 482 82 516
rect 48 410 82 444
rect 48 338 82 372
rect 48 266 82 300
rect 48 194 82 228
rect 454 1058 488 1092
rect 454 986 488 1020
rect 454 914 488 948
rect 454 842 488 876
rect 454 770 488 804
rect 454 698 488 732
rect 454 626 488 660
rect 454 554 488 588
rect 454 482 488 516
rect 454 410 488 444
rect 454 338 488 372
rect 454 266 488 300
rect 454 194 488 228
rect 179 20 213 54
rect 251 20 285 54
rect 323 20 357 54
<< obsli1 >>
rect 159 98 193 1116
rect 251 98 285 1116
rect 343 98 377 1116
<< metal1 >>
rect 167 1194 369 1214
rect 167 1160 179 1194
rect 213 1160 251 1194
rect 285 1160 323 1194
rect 357 1160 369 1194
rect 167 1148 369 1160
rect 36 1092 94 1104
rect 36 1058 48 1092
rect 82 1058 94 1092
rect 36 1020 94 1058
rect 36 986 48 1020
rect 82 986 94 1020
rect 36 948 94 986
rect 36 914 48 948
rect 82 914 94 948
rect 36 876 94 914
rect 36 842 48 876
rect 82 842 94 876
rect 36 804 94 842
rect 36 770 48 804
rect 82 770 94 804
rect 36 732 94 770
rect 36 698 48 732
rect 82 698 94 732
rect 36 660 94 698
rect 36 626 48 660
rect 82 626 94 660
rect 36 588 94 626
rect 36 554 48 588
rect 82 554 94 588
rect 36 516 94 554
rect 36 482 48 516
rect 82 482 94 516
rect 36 444 94 482
rect 36 410 48 444
rect 82 410 94 444
rect 36 372 94 410
rect 36 338 48 372
rect 82 338 94 372
rect 36 300 94 338
rect 36 266 48 300
rect 82 266 94 300
rect 36 228 94 266
rect 36 194 48 228
rect 82 194 94 228
rect 36 110 94 194
rect 442 1092 500 1104
rect 442 1058 454 1092
rect 488 1058 500 1092
rect 442 1020 500 1058
rect 442 986 454 1020
rect 488 986 500 1020
rect 442 948 500 986
rect 442 914 454 948
rect 488 914 500 948
rect 442 876 500 914
rect 442 842 454 876
rect 488 842 500 876
rect 442 804 500 842
rect 442 770 454 804
rect 488 770 500 804
rect 442 732 500 770
rect 442 698 454 732
rect 488 698 500 732
rect 442 660 500 698
rect 442 626 454 660
rect 488 626 500 660
rect 442 588 500 626
rect 442 554 454 588
rect 488 554 500 588
rect 442 516 500 554
rect 442 482 454 516
rect 488 482 500 516
rect 442 444 500 482
rect 442 410 454 444
rect 488 410 500 444
rect 442 372 500 410
rect 442 338 454 372
rect 488 338 500 372
rect 442 300 500 338
rect 442 266 454 300
rect 488 266 500 300
rect 442 228 500 266
rect 442 194 454 228
rect 488 194 500 228
rect 442 110 500 194
rect 167 54 369 66
rect 167 20 179 54
rect 213 20 251 54
rect 285 20 323 54
rect 357 20 369 54
rect 167 0 369 20
<< obsm1 >>
rect 150 110 202 1104
rect 242 110 294 1104
rect 334 110 386 1104
<< metal2 >>
rect 10 632 526 1104
rect 10 110 526 582
<< labels >>
rlabel viali s 454 1058 488 1092 6 BULK
port 1 nsew
rlabel viali s 454 986 488 1020 6 BULK
port 1 nsew
rlabel viali s 454 914 488 948 6 BULK
port 1 nsew
rlabel viali s 454 842 488 876 6 BULK
port 1 nsew
rlabel viali s 454 770 488 804 6 BULK
port 1 nsew
rlabel viali s 454 698 488 732 6 BULK
port 1 nsew
rlabel viali s 454 626 488 660 6 BULK
port 1 nsew
rlabel viali s 454 554 488 588 6 BULK
port 1 nsew
rlabel viali s 454 482 488 516 6 BULK
port 1 nsew
rlabel viali s 454 410 488 444 6 BULK
port 1 nsew
rlabel viali s 454 338 488 372 6 BULK
port 1 nsew
rlabel viali s 454 266 488 300 6 BULK
port 1 nsew
rlabel viali s 454 194 488 228 6 BULK
port 1 nsew
rlabel viali s 48 1058 82 1092 6 BULK
port 1 nsew
rlabel viali s 48 986 82 1020 6 BULK
port 1 nsew
rlabel viali s 48 914 82 948 6 BULK
port 1 nsew
rlabel viali s 48 842 82 876 6 BULK
port 1 nsew
rlabel viali s 48 770 82 804 6 BULK
port 1 nsew
rlabel viali s 48 698 82 732 6 BULK
port 1 nsew
rlabel viali s 48 626 82 660 6 BULK
port 1 nsew
rlabel viali s 48 554 82 588 6 BULK
port 1 nsew
rlabel viali s 48 482 82 516 6 BULK
port 1 nsew
rlabel viali s 48 410 82 444 6 BULK
port 1 nsew
rlabel viali s 48 338 82 372 6 BULK
port 1 nsew
rlabel viali s 48 266 82 300 6 BULK
port 1 nsew
rlabel viali s 48 194 82 228 6 BULK
port 1 nsew
rlabel locali s 454 122 488 1092 6 BULK
port 1 nsew
rlabel locali s 48 122 82 1092 6 BULK
port 1 nsew
rlabel metal1 s 442 110 500 1104 6 BULK
port 1 nsew
rlabel metal1 s 36 110 94 1104 6 BULK
port 1 nsew
rlabel metal2 s 10 632 526 1104 6 DRAIN
port 2 nsew
rlabel viali s 323 1160 357 1194 6 GATE
port 3 nsew
rlabel viali s 323 20 357 54 6 GATE
port 3 nsew
rlabel viali s 251 1160 285 1194 6 GATE
port 3 nsew
rlabel viali s 251 20 285 54 6 GATE
port 3 nsew
rlabel viali s 179 1160 213 1194 6 GATE
port 3 nsew
rlabel viali s 179 20 213 54 6 GATE
port 3 nsew
rlabel locali s 167 1160 369 1194 6 GATE
port 3 nsew
rlabel locali s 167 20 369 54 6 GATE
port 3 nsew
rlabel metal1 s 167 1148 369 1214 6 GATE
port 3 nsew
rlabel metal1 s 167 0 369 66 6 GATE
port 3 nsew
rlabel metal2 s 10 110 526 582 6 SOURCE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 536 1214
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9315700
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9300240
<< end >>
