magic
tech sky130A
magscale 1 2
timestamp 1746986264
<< pwell >>
rect 77 639 87 652
<< obsli1 >>
rect 101 717 371 733
rect 101 683 111 717
rect 145 683 183 717
rect 217 683 255 717
rect 289 683 327 717
rect 361 683 371 717
rect 101 667 371 683
rect 47 605 81 621
rect 47 533 81 571
rect 47 461 81 499
rect 47 389 81 427
rect 47 317 81 355
rect 47 245 81 283
rect 47 173 81 211
rect 47 101 81 139
rect 47 51 81 67
rect 133 51 167 621
rect 219 605 253 621
rect 219 533 253 571
rect 219 461 253 499
rect 219 389 253 427
rect 219 317 253 355
rect 219 245 253 283
rect 219 173 253 211
rect 219 101 253 139
rect 219 51 253 67
rect 305 51 339 621
rect 391 605 425 621
rect 391 533 425 571
rect 391 461 425 499
rect 391 389 425 427
rect 391 317 425 355
rect 391 245 425 283
rect 391 173 425 211
rect 391 101 425 139
rect 391 51 425 67
<< obsli1c >>
rect 111 683 145 717
rect 183 683 217 717
rect 255 683 289 717
rect 327 683 361 717
rect 47 571 81 605
rect 47 499 81 533
rect 47 427 81 461
rect 47 355 81 389
rect 47 283 81 317
rect 47 211 81 245
rect 47 139 81 173
rect 47 67 81 101
rect 219 571 253 605
rect 219 499 253 533
rect 219 427 253 461
rect 219 355 253 389
rect 219 283 253 317
rect 219 211 253 245
rect 219 139 253 173
rect 219 67 253 101
rect 391 571 425 605
rect 391 499 425 533
rect 391 427 425 461
rect 391 355 425 389
rect 391 283 425 317
rect 391 211 425 245
rect 391 139 425 173
rect 391 67 425 101
<< metal1 >>
rect 99 717 373 729
rect 99 683 111 717
rect 145 683 183 717
rect 217 683 255 717
rect 289 683 327 717
rect 361 683 373 717
rect 99 671 373 683
rect 41 605 87 621
rect 41 571 47 605
rect 81 571 87 605
rect 41 533 87 571
rect 41 499 47 533
rect 81 499 87 533
rect 41 461 87 499
rect 41 427 47 461
rect 81 427 87 461
rect 41 389 87 427
rect 41 355 47 389
rect 81 355 87 389
rect 41 317 87 355
rect 41 283 47 317
rect 81 283 87 317
rect 41 245 87 283
rect 41 211 47 245
rect 81 211 87 245
rect 41 173 87 211
rect 41 139 47 173
rect 81 139 87 173
rect 41 101 87 139
rect 41 67 47 101
rect 81 67 87 101
rect 41 -29 87 67
rect 213 605 259 621
rect 213 571 219 605
rect 253 571 259 605
rect 213 533 259 571
rect 213 499 219 533
rect 253 499 259 533
rect 213 461 259 499
rect 213 427 219 461
rect 253 427 259 461
rect 213 389 259 427
rect 213 355 219 389
rect 253 355 259 389
rect 213 317 259 355
rect 213 283 219 317
rect 253 283 259 317
rect 213 245 259 283
rect 213 211 219 245
rect 253 211 259 245
rect 213 173 259 211
rect 213 139 219 173
rect 253 139 259 173
rect 213 101 259 139
rect 213 67 219 101
rect 253 67 259 101
rect 213 -29 259 67
rect 385 605 431 621
rect 385 571 391 605
rect 425 571 431 605
rect 385 533 431 571
rect 385 499 391 533
rect 425 499 431 533
rect 385 461 431 499
rect 385 427 391 461
rect 425 427 431 461
rect 385 389 431 427
rect 385 355 391 389
rect 425 355 431 389
rect 385 317 431 355
rect 385 283 391 317
rect 425 283 431 317
rect 385 245 431 283
rect 385 211 391 245
rect 425 211 431 245
rect 385 173 431 211
rect 385 139 391 173
rect 425 139 431 173
rect 385 101 431 139
rect 385 67 391 101
rect 425 67 431 101
rect 385 -29 431 67
rect 41 -89 431 -29
<< obsm1 >>
rect 124 51 176 621
rect 296 51 348 621
<< obsm2 >>
rect 117 473 183 627
rect 289 473 355 627
<< metal3 >>
rect 117 561 355 627
rect 117 473 183 561
rect 289 473 355 561
<< labels >>
rlabel metal3 s 289 473 355 561 6 DRAIN
port 1 nsew
rlabel metal3 s 117 561 355 627 6 DRAIN
port 1 nsew
rlabel metal3 s 117 473 183 561 6 DRAIN
port 1 nsew
rlabel metal1 s 99 671 373 729 6 GATE
port 2 nsew
rlabel metal1 s 385 -29 431 621 6 SOURCE
port 3 nsew
rlabel metal1 s 213 -29 259 621 6 SOURCE
port 3 nsew
rlabel metal1 s 41 -29 87 621 6 SOURCE
port 3 nsew
rlabel metal1 s 41 -89 431 -29 8 SOURCE
port 3 nsew
rlabel pwell s 77 639 87 652 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 400 822
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10506148
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10495342
string device primitive
<< end >>
